magic
tech sky130A
magscale 1 2
timestamp 1698702074
<< pwell >>
rect -4849 -5082 4849 5082
<< psubdiff >>
rect -4813 5012 -4717 5046
rect 4717 5012 4813 5046
rect -4813 4950 -4779 5012
rect 4779 4950 4813 5012
rect -4813 -5012 -4779 -4950
rect 4779 -5012 4813 -4950
rect -4813 -5046 -4717 -5012
rect 4717 -5046 4813 -5012
<< psubdiffcont >>
rect -4717 5012 4717 5046
rect -4813 -4950 -4779 4950
rect 4779 -4950 4813 4950
rect -4717 -5046 4717 -5012
<< xpolycontact >>
rect -4683 4484 -4613 4916
rect -4683 -4916 -4613 -4484
rect -4517 4484 -4447 4916
rect -4517 -4916 -4447 -4484
rect -4351 4484 -4281 4916
rect -4351 -4916 -4281 -4484
rect -4185 4484 -4115 4916
rect -4185 -4916 -4115 -4484
rect -4019 4484 -3949 4916
rect -4019 -4916 -3949 -4484
rect -3853 4484 -3783 4916
rect -3853 -4916 -3783 -4484
rect -3687 4484 -3617 4916
rect -3687 -4916 -3617 -4484
rect -3521 4484 -3451 4916
rect -3521 -4916 -3451 -4484
rect -3355 4484 -3285 4916
rect -3355 -4916 -3285 -4484
rect -3189 4484 -3119 4916
rect -3189 -4916 -3119 -4484
rect -3023 4484 -2953 4916
rect -3023 -4916 -2953 -4484
rect -2857 4484 -2787 4916
rect -2857 -4916 -2787 -4484
rect -2691 4484 -2621 4916
rect -2691 -4916 -2621 -4484
rect -2525 4484 -2455 4916
rect -2525 -4916 -2455 -4484
rect -2359 4484 -2289 4916
rect -2359 -4916 -2289 -4484
rect -2193 4484 -2123 4916
rect -2193 -4916 -2123 -4484
rect -2027 4484 -1957 4916
rect -2027 -4916 -1957 -4484
rect -1861 4484 -1791 4916
rect -1861 -4916 -1791 -4484
rect -1695 4484 -1625 4916
rect -1695 -4916 -1625 -4484
rect -1529 4484 -1459 4916
rect -1529 -4916 -1459 -4484
rect -1363 4484 -1293 4916
rect -1363 -4916 -1293 -4484
rect -1197 4484 -1127 4916
rect -1197 -4916 -1127 -4484
rect -1031 4484 -961 4916
rect -1031 -4916 -961 -4484
rect -865 4484 -795 4916
rect -865 -4916 -795 -4484
rect -699 4484 -629 4916
rect -699 -4916 -629 -4484
rect -533 4484 -463 4916
rect -533 -4916 -463 -4484
rect -367 4484 -297 4916
rect -367 -4916 -297 -4484
rect -201 4484 -131 4916
rect -201 -4916 -131 -4484
rect -35 4484 35 4916
rect -35 -4916 35 -4484
rect 131 4484 201 4916
rect 131 -4916 201 -4484
rect 297 4484 367 4916
rect 297 -4916 367 -4484
rect 463 4484 533 4916
rect 463 -4916 533 -4484
rect 629 4484 699 4916
rect 629 -4916 699 -4484
rect 795 4484 865 4916
rect 795 -4916 865 -4484
rect 961 4484 1031 4916
rect 961 -4916 1031 -4484
rect 1127 4484 1197 4916
rect 1127 -4916 1197 -4484
rect 1293 4484 1363 4916
rect 1293 -4916 1363 -4484
rect 1459 4484 1529 4916
rect 1459 -4916 1529 -4484
rect 1625 4484 1695 4916
rect 1625 -4916 1695 -4484
rect 1791 4484 1861 4916
rect 1791 -4916 1861 -4484
rect 1957 4484 2027 4916
rect 1957 -4916 2027 -4484
rect 2123 4484 2193 4916
rect 2123 -4916 2193 -4484
rect 2289 4484 2359 4916
rect 2289 -4916 2359 -4484
rect 2455 4484 2525 4916
rect 2455 -4916 2525 -4484
rect 2621 4484 2691 4916
rect 2621 -4916 2691 -4484
rect 2787 4484 2857 4916
rect 2787 -4916 2857 -4484
rect 2953 4484 3023 4916
rect 2953 -4916 3023 -4484
rect 3119 4484 3189 4916
rect 3119 -4916 3189 -4484
rect 3285 4484 3355 4916
rect 3285 -4916 3355 -4484
rect 3451 4484 3521 4916
rect 3451 -4916 3521 -4484
rect 3617 4484 3687 4916
rect 3617 -4916 3687 -4484
rect 3783 4484 3853 4916
rect 3783 -4916 3853 -4484
rect 3949 4484 4019 4916
rect 3949 -4916 4019 -4484
rect 4115 4484 4185 4916
rect 4115 -4916 4185 -4484
rect 4281 4484 4351 4916
rect 4281 -4916 4351 -4484
rect 4447 4484 4517 4916
rect 4447 -4916 4517 -4484
rect 4613 4484 4683 4916
rect 4613 -4916 4683 -4484
<< xpolyres >>
rect -4683 -4484 -4613 4484
rect -4517 -4484 -4447 4484
rect -4351 -4484 -4281 4484
rect -4185 -4484 -4115 4484
rect -4019 -4484 -3949 4484
rect -3853 -4484 -3783 4484
rect -3687 -4484 -3617 4484
rect -3521 -4484 -3451 4484
rect -3355 -4484 -3285 4484
rect -3189 -4484 -3119 4484
rect -3023 -4484 -2953 4484
rect -2857 -4484 -2787 4484
rect -2691 -4484 -2621 4484
rect -2525 -4484 -2455 4484
rect -2359 -4484 -2289 4484
rect -2193 -4484 -2123 4484
rect -2027 -4484 -1957 4484
rect -1861 -4484 -1791 4484
rect -1695 -4484 -1625 4484
rect -1529 -4484 -1459 4484
rect -1363 -4484 -1293 4484
rect -1197 -4484 -1127 4484
rect -1031 -4484 -961 4484
rect -865 -4484 -795 4484
rect -699 -4484 -629 4484
rect -533 -4484 -463 4484
rect -367 -4484 -297 4484
rect -201 -4484 -131 4484
rect -35 -4484 35 4484
rect 131 -4484 201 4484
rect 297 -4484 367 4484
rect 463 -4484 533 4484
rect 629 -4484 699 4484
rect 795 -4484 865 4484
rect 961 -4484 1031 4484
rect 1127 -4484 1197 4484
rect 1293 -4484 1363 4484
rect 1459 -4484 1529 4484
rect 1625 -4484 1695 4484
rect 1791 -4484 1861 4484
rect 1957 -4484 2027 4484
rect 2123 -4484 2193 4484
rect 2289 -4484 2359 4484
rect 2455 -4484 2525 4484
rect 2621 -4484 2691 4484
rect 2787 -4484 2857 4484
rect 2953 -4484 3023 4484
rect 3119 -4484 3189 4484
rect 3285 -4484 3355 4484
rect 3451 -4484 3521 4484
rect 3617 -4484 3687 4484
rect 3783 -4484 3853 4484
rect 3949 -4484 4019 4484
rect 4115 -4484 4185 4484
rect 4281 -4484 4351 4484
rect 4447 -4484 4517 4484
rect 4613 -4484 4683 4484
<< locali >>
rect -4813 5012 -4717 5046
rect 4717 5012 4813 5046
rect -4813 4950 -4779 5012
rect 4779 4950 4813 5012
rect -4813 -5012 -4779 -4950
rect 4779 -5012 4813 -4950
rect -4813 -5046 -4717 -5012
rect 4717 -5046 4813 -5012
<< viali >>
rect -4667 4501 -4629 4898
rect -4501 4501 -4463 4898
rect -4335 4501 -4297 4898
rect -4169 4501 -4131 4898
rect -4003 4501 -3965 4898
rect -3837 4501 -3799 4898
rect -3671 4501 -3633 4898
rect -3505 4501 -3467 4898
rect -3339 4501 -3301 4898
rect -3173 4501 -3135 4898
rect -3007 4501 -2969 4898
rect -2841 4501 -2803 4898
rect -2675 4501 -2637 4898
rect -2509 4501 -2471 4898
rect -2343 4501 -2305 4898
rect -2177 4501 -2139 4898
rect -2011 4501 -1973 4898
rect -1845 4501 -1807 4898
rect -1679 4501 -1641 4898
rect -1513 4501 -1475 4898
rect -1347 4501 -1309 4898
rect -1181 4501 -1143 4898
rect -1015 4501 -977 4898
rect -849 4501 -811 4898
rect -683 4501 -645 4898
rect -517 4501 -479 4898
rect -351 4501 -313 4898
rect -185 4501 -147 4898
rect -19 4501 19 4898
rect 147 4501 185 4898
rect 313 4501 351 4898
rect 479 4501 517 4898
rect 645 4501 683 4898
rect 811 4501 849 4898
rect 977 4501 1015 4898
rect 1143 4501 1181 4898
rect 1309 4501 1347 4898
rect 1475 4501 1513 4898
rect 1641 4501 1679 4898
rect 1807 4501 1845 4898
rect 1973 4501 2011 4898
rect 2139 4501 2177 4898
rect 2305 4501 2343 4898
rect 2471 4501 2509 4898
rect 2637 4501 2675 4898
rect 2803 4501 2841 4898
rect 2969 4501 3007 4898
rect 3135 4501 3173 4898
rect 3301 4501 3339 4898
rect 3467 4501 3505 4898
rect 3633 4501 3671 4898
rect 3799 4501 3837 4898
rect 3965 4501 4003 4898
rect 4131 4501 4169 4898
rect 4297 4501 4335 4898
rect 4463 4501 4501 4898
rect 4629 4501 4667 4898
rect -4667 -4898 -4629 -4501
rect -4501 -4898 -4463 -4501
rect -4335 -4898 -4297 -4501
rect -4169 -4898 -4131 -4501
rect -4003 -4898 -3965 -4501
rect -3837 -4898 -3799 -4501
rect -3671 -4898 -3633 -4501
rect -3505 -4898 -3467 -4501
rect -3339 -4898 -3301 -4501
rect -3173 -4898 -3135 -4501
rect -3007 -4898 -2969 -4501
rect -2841 -4898 -2803 -4501
rect -2675 -4898 -2637 -4501
rect -2509 -4898 -2471 -4501
rect -2343 -4898 -2305 -4501
rect -2177 -4898 -2139 -4501
rect -2011 -4898 -1973 -4501
rect -1845 -4898 -1807 -4501
rect -1679 -4898 -1641 -4501
rect -1513 -4898 -1475 -4501
rect -1347 -4898 -1309 -4501
rect -1181 -4898 -1143 -4501
rect -1015 -4898 -977 -4501
rect -849 -4898 -811 -4501
rect -683 -4898 -645 -4501
rect -517 -4898 -479 -4501
rect -351 -4898 -313 -4501
rect -185 -4898 -147 -4501
rect -19 -4898 19 -4501
rect 147 -4898 185 -4501
rect 313 -4898 351 -4501
rect 479 -4898 517 -4501
rect 645 -4898 683 -4501
rect 811 -4898 849 -4501
rect 977 -4898 1015 -4501
rect 1143 -4898 1181 -4501
rect 1309 -4898 1347 -4501
rect 1475 -4898 1513 -4501
rect 1641 -4898 1679 -4501
rect 1807 -4898 1845 -4501
rect 1973 -4898 2011 -4501
rect 2139 -4898 2177 -4501
rect 2305 -4898 2343 -4501
rect 2471 -4898 2509 -4501
rect 2637 -4898 2675 -4501
rect 2803 -4898 2841 -4501
rect 2969 -4898 3007 -4501
rect 3135 -4898 3173 -4501
rect 3301 -4898 3339 -4501
rect 3467 -4898 3505 -4501
rect 3633 -4898 3671 -4501
rect 3799 -4898 3837 -4501
rect 3965 -4898 4003 -4501
rect 4131 -4898 4169 -4501
rect 4297 -4898 4335 -4501
rect 4463 -4898 4501 -4501
rect 4629 -4898 4667 -4501
<< metal1 >>
rect -4673 4898 -4623 4910
rect -4673 4501 -4667 4898
rect -4629 4501 -4623 4898
rect -4673 4489 -4623 4501
rect -4507 4898 -4457 4910
rect -4507 4501 -4501 4898
rect -4463 4501 -4457 4898
rect -4507 4489 -4457 4501
rect -4341 4898 -4291 4910
rect -4341 4501 -4335 4898
rect -4297 4501 -4291 4898
rect -4341 4489 -4291 4501
rect -4175 4898 -4125 4910
rect -4175 4501 -4169 4898
rect -4131 4501 -4125 4898
rect -4175 4489 -4125 4501
rect -4009 4898 -3959 4910
rect -4009 4501 -4003 4898
rect -3965 4501 -3959 4898
rect -4009 4489 -3959 4501
rect -3843 4898 -3793 4910
rect -3843 4501 -3837 4898
rect -3799 4501 -3793 4898
rect -3843 4489 -3793 4501
rect -3677 4898 -3627 4910
rect -3677 4501 -3671 4898
rect -3633 4501 -3627 4898
rect -3677 4489 -3627 4501
rect -3511 4898 -3461 4910
rect -3511 4501 -3505 4898
rect -3467 4501 -3461 4898
rect -3511 4489 -3461 4501
rect -3345 4898 -3295 4910
rect -3345 4501 -3339 4898
rect -3301 4501 -3295 4898
rect -3345 4489 -3295 4501
rect -3179 4898 -3129 4910
rect -3179 4501 -3173 4898
rect -3135 4501 -3129 4898
rect -3179 4489 -3129 4501
rect -3013 4898 -2963 4910
rect -3013 4501 -3007 4898
rect -2969 4501 -2963 4898
rect -3013 4489 -2963 4501
rect -2847 4898 -2797 4910
rect -2847 4501 -2841 4898
rect -2803 4501 -2797 4898
rect -2847 4489 -2797 4501
rect -2681 4898 -2631 4910
rect -2681 4501 -2675 4898
rect -2637 4501 -2631 4898
rect -2681 4489 -2631 4501
rect -2515 4898 -2465 4910
rect -2515 4501 -2509 4898
rect -2471 4501 -2465 4898
rect -2515 4489 -2465 4501
rect -2349 4898 -2299 4910
rect -2349 4501 -2343 4898
rect -2305 4501 -2299 4898
rect -2349 4489 -2299 4501
rect -2183 4898 -2133 4910
rect -2183 4501 -2177 4898
rect -2139 4501 -2133 4898
rect -2183 4489 -2133 4501
rect -2017 4898 -1967 4910
rect -2017 4501 -2011 4898
rect -1973 4501 -1967 4898
rect -2017 4489 -1967 4501
rect -1851 4898 -1801 4910
rect -1851 4501 -1845 4898
rect -1807 4501 -1801 4898
rect -1851 4489 -1801 4501
rect -1685 4898 -1635 4910
rect -1685 4501 -1679 4898
rect -1641 4501 -1635 4898
rect -1685 4489 -1635 4501
rect -1519 4898 -1469 4910
rect -1519 4501 -1513 4898
rect -1475 4501 -1469 4898
rect -1519 4489 -1469 4501
rect -1353 4898 -1303 4910
rect -1353 4501 -1347 4898
rect -1309 4501 -1303 4898
rect -1353 4489 -1303 4501
rect -1187 4898 -1137 4910
rect -1187 4501 -1181 4898
rect -1143 4501 -1137 4898
rect -1187 4489 -1137 4501
rect -1021 4898 -971 4910
rect -1021 4501 -1015 4898
rect -977 4501 -971 4898
rect -1021 4489 -971 4501
rect -855 4898 -805 4910
rect -855 4501 -849 4898
rect -811 4501 -805 4898
rect -855 4489 -805 4501
rect -689 4898 -639 4910
rect -689 4501 -683 4898
rect -645 4501 -639 4898
rect -689 4489 -639 4501
rect -523 4898 -473 4910
rect -523 4501 -517 4898
rect -479 4501 -473 4898
rect -523 4489 -473 4501
rect -357 4898 -307 4910
rect -357 4501 -351 4898
rect -313 4501 -307 4898
rect -357 4489 -307 4501
rect -191 4898 -141 4910
rect -191 4501 -185 4898
rect -147 4501 -141 4898
rect -191 4489 -141 4501
rect -25 4898 25 4910
rect -25 4501 -19 4898
rect 19 4501 25 4898
rect -25 4489 25 4501
rect 141 4898 191 4910
rect 141 4501 147 4898
rect 185 4501 191 4898
rect 141 4489 191 4501
rect 307 4898 357 4910
rect 307 4501 313 4898
rect 351 4501 357 4898
rect 307 4489 357 4501
rect 473 4898 523 4910
rect 473 4501 479 4898
rect 517 4501 523 4898
rect 473 4489 523 4501
rect 639 4898 689 4910
rect 639 4501 645 4898
rect 683 4501 689 4898
rect 639 4489 689 4501
rect 805 4898 855 4910
rect 805 4501 811 4898
rect 849 4501 855 4898
rect 805 4489 855 4501
rect 971 4898 1021 4910
rect 971 4501 977 4898
rect 1015 4501 1021 4898
rect 971 4489 1021 4501
rect 1137 4898 1187 4910
rect 1137 4501 1143 4898
rect 1181 4501 1187 4898
rect 1137 4489 1187 4501
rect 1303 4898 1353 4910
rect 1303 4501 1309 4898
rect 1347 4501 1353 4898
rect 1303 4489 1353 4501
rect 1469 4898 1519 4910
rect 1469 4501 1475 4898
rect 1513 4501 1519 4898
rect 1469 4489 1519 4501
rect 1635 4898 1685 4910
rect 1635 4501 1641 4898
rect 1679 4501 1685 4898
rect 1635 4489 1685 4501
rect 1801 4898 1851 4910
rect 1801 4501 1807 4898
rect 1845 4501 1851 4898
rect 1801 4489 1851 4501
rect 1967 4898 2017 4910
rect 1967 4501 1973 4898
rect 2011 4501 2017 4898
rect 1967 4489 2017 4501
rect 2133 4898 2183 4910
rect 2133 4501 2139 4898
rect 2177 4501 2183 4898
rect 2133 4489 2183 4501
rect 2299 4898 2349 4910
rect 2299 4501 2305 4898
rect 2343 4501 2349 4898
rect 2299 4489 2349 4501
rect 2465 4898 2515 4910
rect 2465 4501 2471 4898
rect 2509 4501 2515 4898
rect 2465 4489 2515 4501
rect 2631 4898 2681 4910
rect 2631 4501 2637 4898
rect 2675 4501 2681 4898
rect 2631 4489 2681 4501
rect 2797 4898 2847 4910
rect 2797 4501 2803 4898
rect 2841 4501 2847 4898
rect 2797 4489 2847 4501
rect 2963 4898 3013 4910
rect 2963 4501 2969 4898
rect 3007 4501 3013 4898
rect 2963 4489 3013 4501
rect 3129 4898 3179 4910
rect 3129 4501 3135 4898
rect 3173 4501 3179 4898
rect 3129 4489 3179 4501
rect 3295 4898 3345 4910
rect 3295 4501 3301 4898
rect 3339 4501 3345 4898
rect 3295 4489 3345 4501
rect 3461 4898 3511 4910
rect 3461 4501 3467 4898
rect 3505 4501 3511 4898
rect 3461 4489 3511 4501
rect 3627 4898 3677 4910
rect 3627 4501 3633 4898
rect 3671 4501 3677 4898
rect 3627 4489 3677 4501
rect 3793 4898 3843 4910
rect 3793 4501 3799 4898
rect 3837 4501 3843 4898
rect 3793 4489 3843 4501
rect 3959 4898 4009 4910
rect 3959 4501 3965 4898
rect 4003 4501 4009 4898
rect 3959 4489 4009 4501
rect 4125 4898 4175 4910
rect 4125 4501 4131 4898
rect 4169 4501 4175 4898
rect 4125 4489 4175 4501
rect 4291 4898 4341 4910
rect 4291 4501 4297 4898
rect 4335 4501 4341 4898
rect 4291 4489 4341 4501
rect 4457 4898 4507 4910
rect 4457 4501 4463 4898
rect 4501 4501 4507 4898
rect 4457 4489 4507 4501
rect 4623 4898 4673 4910
rect 4623 4501 4629 4898
rect 4667 4501 4673 4898
rect 4623 4489 4673 4501
rect -4673 -4501 -4623 -4489
rect -4673 -4898 -4667 -4501
rect -4629 -4898 -4623 -4501
rect -4673 -4910 -4623 -4898
rect -4507 -4501 -4457 -4489
rect -4507 -4898 -4501 -4501
rect -4463 -4898 -4457 -4501
rect -4507 -4910 -4457 -4898
rect -4341 -4501 -4291 -4489
rect -4341 -4898 -4335 -4501
rect -4297 -4898 -4291 -4501
rect -4341 -4910 -4291 -4898
rect -4175 -4501 -4125 -4489
rect -4175 -4898 -4169 -4501
rect -4131 -4898 -4125 -4501
rect -4175 -4910 -4125 -4898
rect -4009 -4501 -3959 -4489
rect -4009 -4898 -4003 -4501
rect -3965 -4898 -3959 -4501
rect -4009 -4910 -3959 -4898
rect -3843 -4501 -3793 -4489
rect -3843 -4898 -3837 -4501
rect -3799 -4898 -3793 -4501
rect -3843 -4910 -3793 -4898
rect -3677 -4501 -3627 -4489
rect -3677 -4898 -3671 -4501
rect -3633 -4898 -3627 -4501
rect -3677 -4910 -3627 -4898
rect -3511 -4501 -3461 -4489
rect -3511 -4898 -3505 -4501
rect -3467 -4898 -3461 -4501
rect -3511 -4910 -3461 -4898
rect -3345 -4501 -3295 -4489
rect -3345 -4898 -3339 -4501
rect -3301 -4898 -3295 -4501
rect -3345 -4910 -3295 -4898
rect -3179 -4501 -3129 -4489
rect -3179 -4898 -3173 -4501
rect -3135 -4898 -3129 -4501
rect -3179 -4910 -3129 -4898
rect -3013 -4501 -2963 -4489
rect -3013 -4898 -3007 -4501
rect -2969 -4898 -2963 -4501
rect -3013 -4910 -2963 -4898
rect -2847 -4501 -2797 -4489
rect -2847 -4898 -2841 -4501
rect -2803 -4898 -2797 -4501
rect -2847 -4910 -2797 -4898
rect -2681 -4501 -2631 -4489
rect -2681 -4898 -2675 -4501
rect -2637 -4898 -2631 -4501
rect -2681 -4910 -2631 -4898
rect -2515 -4501 -2465 -4489
rect -2515 -4898 -2509 -4501
rect -2471 -4898 -2465 -4501
rect -2515 -4910 -2465 -4898
rect -2349 -4501 -2299 -4489
rect -2349 -4898 -2343 -4501
rect -2305 -4898 -2299 -4501
rect -2349 -4910 -2299 -4898
rect -2183 -4501 -2133 -4489
rect -2183 -4898 -2177 -4501
rect -2139 -4898 -2133 -4501
rect -2183 -4910 -2133 -4898
rect -2017 -4501 -1967 -4489
rect -2017 -4898 -2011 -4501
rect -1973 -4898 -1967 -4501
rect -2017 -4910 -1967 -4898
rect -1851 -4501 -1801 -4489
rect -1851 -4898 -1845 -4501
rect -1807 -4898 -1801 -4501
rect -1851 -4910 -1801 -4898
rect -1685 -4501 -1635 -4489
rect -1685 -4898 -1679 -4501
rect -1641 -4898 -1635 -4501
rect -1685 -4910 -1635 -4898
rect -1519 -4501 -1469 -4489
rect -1519 -4898 -1513 -4501
rect -1475 -4898 -1469 -4501
rect -1519 -4910 -1469 -4898
rect -1353 -4501 -1303 -4489
rect -1353 -4898 -1347 -4501
rect -1309 -4898 -1303 -4501
rect -1353 -4910 -1303 -4898
rect -1187 -4501 -1137 -4489
rect -1187 -4898 -1181 -4501
rect -1143 -4898 -1137 -4501
rect -1187 -4910 -1137 -4898
rect -1021 -4501 -971 -4489
rect -1021 -4898 -1015 -4501
rect -977 -4898 -971 -4501
rect -1021 -4910 -971 -4898
rect -855 -4501 -805 -4489
rect -855 -4898 -849 -4501
rect -811 -4898 -805 -4501
rect -855 -4910 -805 -4898
rect -689 -4501 -639 -4489
rect -689 -4898 -683 -4501
rect -645 -4898 -639 -4501
rect -689 -4910 -639 -4898
rect -523 -4501 -473 -4489
rect -523 -4898 -517 -4501
rect -479 -4898 -473 -4501
rect -523 -4910 -473 -4898
rect -357 -4501 -307 -4489
rect -357 -4898 -351 -4501
rect -313 -4898 -307 -4501
rect -357 -4910 -307 -4898
rect -191 -4501 -141 -4489
rect -191 -4898 -185 -4501
rect -147 -4898 -141 -4501
rect -191 -4910 -141 -4898
rect -25 -4501 25 -4489
rect -25 -4898 -19 -4501
rect 19 -4898 25 -4501
rect -25 -4910 25 -4898
rect 141 -4501 191 -4489
rect 141 -4898 147 -4501
rect 185 -4898 191 -4501
rect 141 -4910 191 -4898
rect 307 -4501 357 -4489
rect 307 -4898 313 -4501
rect 351 -4898 357 -4501
rect 307 -4910 357 -4898
rect 473 -4501 523 -4489
rect 473 -4898 479 -4501
rect 517 -4898 523 -4501
rect 473 -4910 523 -4898
rect 639 -4501 689 -4489
rect 639 -4898 645 -4501
rect 683 -4898 689 -4501
rect 639 -4910 689 -4898
rect 805 -4501 855 -4489
rect 805 -4898 811 -4501
rect 849 -4898 855 -4501
rect 805 -4910 855 -4898
rect 971 -4501 1021 -4489
rect 971 -4898 977 -4501
rect 1015 -4898 1021 -4501
rect 971 -4910 1021 -4898
rect 1137 -4501 1187 -4489
rect 1137 -4898 1143 -4501
rect 1181 -4898 1187 -4501
rect 1137 -4910 1187 -4898
rect 1303 -4501 1353 -4489
rect 1303 -4898 1309 -4501
rect 1347 -4898 1353 -4501
rect 1303 -4910 1353 -4898
rect 1469 -4501 1519 -4489
rect 1469 -4898 1475 -4501
rect 1513 -4898 1519 -4501
rect 1469 -4910 1519 -4898
rect 1635 -4501 1685 -4489
rect 1635 -4898 1641 -4501
rect 1679 -4898 1685 -4501
rect 1635 -4910 1685 -4898
rect 1801 -4501 1851 -4489
rect 1801 -4898 1807 -4501
rect 1845 -4898 1851 -4501
rect 1801 -4910 1851 -4898
rect 1967 -4501 2017 -4489
rect 1967 -4898 1973 -4501
rect 2011 -4898 2017 -4501
rect 1967 -4910 2017 -4898
rect 2133 -4501 2183 -4489
rect 2133 -4898 2139 -4501
rect 2177 -4898 2183 -4501
rect 2133 -4910 2183 -4898
rect 2299 -4501 2349 -4489
rect 2299 -4898 2305 -4501
rect 2343 -4898 2349 -4501
rect 2299 -4910 2349 -4898
rect 2465 -4501 2515 -4489
rect 2465 -4898 2471 -4501
rect 2509 -4898 2515 -4501
rect 2465 -4910 2515 -4898
rect 2631 -4501 2681 -4489
rect 2631 -4898 2637 -4501
rect 2675 -4898 2681 -4501
rect 2631 -4910 2681 -4898
rect 2797 -4501 2847 -4489
rect 2797 -4898 2803 -4501
rect 2841 -4898 2847 -4501
rect 2797 -4910 2847 -4898
rect 2963 -4501 3013 -4489
rect 2963 -4898 2969 -4501
rect 3007 -4898 3013 -4501
rect 2963 -4910 3013 -4898
rect 3129 -4501 3179 -4489
rect 3129 -4898 3135 -4501
rect 3173 -4898 3179 -4501
rect 3129 -4910 3179 -4898
rect 3295 -4501 3345 -4489
rect 3295 -4898 3301 -4501
rect 3339 -4898 3345 -4501
rect 3295 -4910 3345 -4898
rect 3461 -4501 3511 -4489
rect 3461 -4898 3467 -4501
rect 3505 -4898 3511 -4501
rect 3461 -4910 3511 -4898
rect 3627 -4501 3677 -4489
rect 3627 -4898 3633 -4501
rect 3671 -4898 3677 -4501
rect 3627 -4910 3677 -4898
rect 3793 -4501 3843 -4489
rect 3793 -4898 3799 -4501
rect 3837 -4898 3843 -4501
rect 3793 -4910 3843 -4898
rect 3959 -4501 4009 -4489
rect 3959 -4898 3965 -4501
rect 4003 -4898 4009 -4501
rect 3959 -4910 4009 -4898
rect 4125 -4501 4175 -4489
rect 4125 -4898 4131 -4501
rect 4169 -4898 4175 -4501
rect 4125 -4910 4175 -4898
rect 4291 -4501 4341 -4489
rect 4291 -4898 4297 -4501
rect 4335 -4898 4341 -4501
rect 4291 -4910 4341 -4898
rect 4457 -4501 4507 -4489
rect 4457 -4898 4463 -4501
rect 4501 -4898 4507 -4501
rect 4457 -4910 4507 -4898
rect 4623 -4501 4673 -4489
rect 4623 -4898 4629 -4501
rect 4667 -4898 4673 -4501
rect 4623 -4910 4673 -4898
<< properties >>
string FIXED_BBOX -4796 -5029 4796 5029
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 45.0 m 1 nx 57 wmin 0.350 lmin 0.50 rho 2000 val 258.218k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
