magic
tech sky130A
magscale 1 2
timestamp 1698702074
<< pwell >>
rect -1695 -5082 1695 5082
<< psubdiff >>
rect -1659 5012 -1563 5046
rect 1563 5012 1659 5046
rect -1659 4950 -1625 5012
rect 1625 4950 1659 5012
rect -1659 -5012 -1625 -4950
rect 1625 -5012 1659 -4950
rect -1659 -5046 -1563 -5012
rect 1563 -5046 1659 -5012
<< psubdiffcont >>
rect -1563 5012 1563 5046
rect -1659 -4950 -1625 4950
rect 1625 -4950 1659 4950
rect -1563 -5046 1563 -5012
<< xpolycontact >>
rect -1529 4484 -1459 4916
rect -1529 -4916 -1459 -4484
rect -1363 4484 -1293 4916
rect -1363 -4916 -1293 -4484
rect -1197 4484 -1127 4916
rect -1197 -4916 -1127 -4484
rect -1031 4484 -961 4916
rect -1031 -4916 -961 -4484
rect -865 4484 -795 4916
rect -865 -4916 -795 -4484
rect -699 4484 -629 4916
rect -699 -4916 -629 -4484
rect -533 4484 -463 4916
rect -533 -4916 -463 -4484
rect -367 4484 -297 4916
rect -367 -4916 -297 -4484
rect -201 4484 -131 4916
rect -201 -4916 -131 -4484
rect -35 4484 35 4916
rect -35 -4916 35 -4484
rect 131 4484 201 4916
rect 131 -4916 201 -4484
rect 297 4484 367 4916
rect 297 -4916 367 -4484
rect 463 4484 533 4916
rect 463 -4916 533 -4484
rect 629 4484 699 4916
rect 629 -4916 699 -4484
rect 795 4484 865 4916
rect 795 -4916 865 -4484
rect 961 4484 1031 4916
rect 961 -4916 1031 -4484
rect 1127 4484 1197 4916
rect 1127 -4916 1197 -4484
rect 1293 4484 1363 4916
rect 1293 -4916 1363 -4484
rect 1459 4484 1529 4916
rect 1459 -4916 1529 -4484
<< xpolyres >>
rect -1529 -4484 -1459 4484
rect -1363 -4484 -1293 4484
rect -1197 -4484 -1127 4484
rect -1031 -4484 -961 4484
rect -865 -4484 -795 4484
rect -699 -4484 -629 4484
rect -533 -4484 -463 4484
rect -367 -4484 -297 4484
rect -201 -4484 -131 4484
rect -35 -4484 35 4484
rect 131 -4484 201 4484
rect 297 -4484 367 4484
rect 463 -4484 533 4484
rect 629 -4484 699 4484
rect 795 -4484 865 4484
rect 961 -4484 1031 4484
rect 1127 -4484 1197 4484
rect 1293 -4484 1363 4484
rect 1459 -4484 1529 4484
<< locali >>
rect -1659 5012 -1563 5046
rect 1563 5012 1659 5046
rect -1659 4950 -1625 5012
rect 1625 4950 1659 5012
rect -1659 -5012 -1625 -4950
rect 1625 -5012 1659 -4950
rect -1659 -5046 -1563 -5012
rect 1563 -5046 1659 -5012
<< viali >>
rect -1513 4501 -1475 4898
rect -1347 4501 -1309 4898
rect -1181 4501 -1143 4898
rect -1015 4501 -977 4898
rect -849 4501 -811 4898
rect -683 4501 -645 4898
rect -517 4501 -479 4898
rect -351 4501 -313 4898
rect -185 4501 -147 4898
rect -19 4501 19 4898
rect 147 4501 185 4898
rect 313 4501 351 4898
rect 479 4501 517 4898
rect 645 4501 683 4898
rect 811 4501 849 4898
rect 977 4501 1015 4898
rect 1143 4501 1181 4898
rect 1309 4501 1347 4898
rect 1475 4501 1513 4898
rect -1513 -4898 -1475 -4501
rect -1347 -4898 -1309 -4501
rect -1181 -4898 -1143 -4501
rect -1015 -4898 -977 -4501
rect -849 -4898 -811 -4501
rect -683 -4898 -645 -4501
rect -517 -4898 -479 -4501
rect -351 -4898 -313 -4501
rect -185 -4898 -147 -4501
rect -19 -4898 19 -4501
rect 147 -4898 185 -4501
rect 313 -4898 351 -4501
rect 479 -4898 517 -4501
rect 645 -4898 683 -4501
rect 811 -4898 849 -4501
rect 977 -4898 1015 -4501
rect 1143 -4898 1181 -4501
rect 1309 -4898 1347 -4501
rect 1475 -4898 1513 -4501
<< metal1 >>
rect -1519 4898 -1469 4910
rect -1519 4501 -1513 4898
rect -1475 4501 -1469 4898
rect -1519 4489 -1469 4501
rect -1353 4898 -1303 4910
rect -1353 4501 -1347 4898
rect -1309 4501 -1303 4898
rect -1353 4489 -1303 4501
rect -1187 4898 -1137 4910
rect -1187 4501 -1181 4898
rect -1143 4501 -1137 4898
rect -1187 4489 -1137 4501
rect -1021 4898 -971 4910
rect -1021 4501 -1015 4898
rect -977 4501 -971 4898
rect -1021 4489 -971 4501
rect -855 4898 -805 4910
rect -855 4501 -849 4898
rect -811 4501 -805 4898
rect -855 4489 -805 4501
rect -689 4898 -639 4910
rect -689 4501 -683 4898
rect -645 4501 -639 4898
rect -689 4489 -639 4501
rect -523 4898 -473 4910
rect -523 4501 -517 4898
rect -479 4501 -473 4898
rect -523 4489 -473 4501
rect -357 4898 -307 4910
rect -357 4501 -351 4898
rect -313 4501 -307 4898
rect -357 4489 -307 4501
rect -191 4898 -141 4910
rect -191 4501 -185 4898
rect -147 4501 -141 4898
rect -191 4489 -141 4501
rect -25 4898 25 4910
rect -25 4501 -19 4898
rect 19 4501 25 4898
rect -25 4489 25 4501
rect 141 4898 191 4910
rect 141 4501 147 4898
rect 185 4501 191 4898
rect 141 4489 191 4501
rect 307 4898 357 4910
rect 307 4501 313 4898
rect 351 4501 357 4898
rect 307 4489 357 4501
rect 473 4898 523 4910
rect 473 4501 479 4898
rect 517 4501 523 4898
rect 473 4489 523 4501
rect 639 4898 689 4910
rect 639 4501 645 4898
rect 683 4501 689 4898
rect 639 4489 689 4501
rect 805 4898 855 4910
rect 805 4501 811 4898
rect 849 4501 855 4898
rect 805 4489 855 4501
rect 971 4898 1021 4910
rect 971 4501 977 4898
rect 1015 4501 1021 4898
rect 971 4489 1021 4501
rect 1137 4898 1187 4910
rect 1137 4501 1143 4898
rect 1181 4501 1187 4898
rect 1137 4489 1187 4501
rect 1303 4898 1353 4910
rect 1303 4501 1309 4898
rect 1347 4501 1353 4898
rect 1303 4489 1353 4501
rect 1469 4898 1519 4910
rect 1469 4501 1475 4898
rect 1513 4501 1519 4898
rect 1469 4489 1519 4501
rect -1519 -4501 -1469 -4489
rect -1519 -4898 -1513 -4501
rect -1475 -4898 -1469 -4501
rect -1519 -4910 -1469 -4898
rect -1353 -4501 -1303 -4489
rect -1353 -4898 -1347 -4501
rect -1309 -4898 -1303 -4501
rect -1353 -4910 -1303 -4898
rect -1187 -4501 -1137 -4489
rect -1187 -4898 -1181 -4501
rect -1143 -4898 -1137 -4501
rect -1187 -4910 -1137 -4898
rect -1021 -4501 -971 -4489
rect -1021 -4898 -1015 -4501
rect -977 -4898 -971 -4501
rect -1021 -4910 -971 -4898
rect -855 -4501 -805 -4489
rect -855 -4898 -849 -4501
rect -811 -4898 -805 -4501
rect -855 -4910 -805 -4898
rect -689 -4501 -639 -4489
rect -689 -4898 -683 -4501
rect -645 -4898 -639 -4501
rect -689 -4910 -639 -4898
rect -523 -4501 -473 -4489
rect -523 -4898 -517 -4501
rect -479 -4898 -473 -4501
rect -523 -4910 -473 -4898
rect -357 -4501 -307 -4489
rect -357 -4898 -351 -4501
rect -313 -4898 -307 -4501
rect -357 -4910 -307 -4898
rect -191 -4501 -141 -4489
rect -191 -4898 -185 -4501
rect -147 -4898 -141 -4501
rect -191 -4910 -141 -4898
rect -25 -4501 25 -4489
rect -25 -4898 -19 -4501
rect 19 -4898 25 -4501
rect -25 -4910 25 -4898
rect 141 -4501 191 -4489
rect 141 -4898 147 -4501
rect 185 -4898 191 -4501
rect 141 -4910 191 -4898
rect 307 -4501 357 -4489
rect 307 -4898 313 -4501
rect 351 -4898 357 -4501
rect 307 -4910 357 -4898
rect 473 -4501 523 -4489
rect 473 -4898 479 -4501
rect 517 -4898 523 -4501
rect 473 -4910 523 -4898
rect 639 -4501 689 -4489
rect 639 -4898 645 -4501
rect 683 -4898 689 -4501
rect 639 -4910 689 -4898
rect 805 -4501 855 -4489
rect 805 -4898 811 -4501
rect 849 -4898 855 -4501
rect 805 -4910 855 -4898
rect 971 -4501 1021 -4489
rect 971 -4898 977 -4501
rect 1015 -4898 1021 -4501
rect 971 -4910 1021 -4898
rect 1137 -4501 1187 -4489
rect 1137 -4898 1143 -4501
rect 1181 -4898 1187 -4501
rect 1137 -4910 1187 -4898
rect 1303 -4501 1353 -4489
rect 1303 -4898 1309 -4501
rect 1347 -4898 1353 -4501
rect 1303 -4910 1353 -4898
rect 1469 -4501 1519 -4489
rect 1469 -4898 1475 -4501
rect 1513 -4898 1519 -4501
rect 1469 -4910 1519 -4898
<< properties >>
string FIXED_BBOX -1642 -5029 1642 5029
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 45.0 m 1 nx 19 wmin 0.350 lmin 0.50 rho 2000 val 258.218k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
