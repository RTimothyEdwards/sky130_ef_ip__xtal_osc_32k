magic
tech sky130A
magscale 1 2
timestamp 1698863670
<< dnwell >>
rect 10988 -1960 24802 8744
rect 10988 -6898 23092 -1960
rect 10988 -17594 24802 -6898
<< nwell >>
rect 10878 8538 24912 8854
rect 10878 -17358 11194 8538
rect 24596 -1752 24912 8538
rect 22886 -2068 24912 -1752
rect 17712 -3586 18328 -2978
rect 20792 -3586 20884 -2978
rect 22886 -3000 23202 -2068
rect 17712 -3656 20884 -3586
rect 20792 -4264 20884 -3656
rect 22858 -4346 23202 -3000
rect 24414 -3846 24500 -3278
rect 21632 -4570 23202 -4346
rect 22858 -5907 23202 -4570
rect 22886 -6788 23202 -5907
rect 22886 -7104 24912 -6788
rect 24596 -17358 24912 -7104
rect 10878 -17704 24912 -17358
<< mvnsubdiff >>
rect 10945 8767 24845 8787
rect 10945 8733 11025 8767
rect 24765 8733 24845 8767
rect 10945 8713 24845 8733
rect 10945 8707 11019 8713
rect 10945 -17557 10965 8707
rect 10999 -17557 11019 8707
rect 24771 8707 24845 8713
rect 24771 -1906 24791 8707
rect 24825 -1906 24845 8707
rect 24771 -1925 24845 -1906
rect 23051 -1945 24845 -1925
rect 23051 -1979 23145 -1945
rect 24775 -1979 24845 -1945
rect 23051 -1995 24845 -1979
rect 23051 -6871 23071 -1995
rect 23105 -1999 24845 -1995
rect 23105 -6867 23125 -1999
rect 23105 -6871 24845 -6867
rect 23051 -6887 24845 -6871
rect 23051 -6921 23141 -6887
rect 24755 -6921 24845 -6887
rect 23051 -6941 24845 -6921
rect 10945 -17563 11019 -17557
rect 24771 -6956 24845 -6941
rect 24771 -17554 24791 -6956
rect 24825 -17554 24845 -6956
rect 24771 -17563 24845 -17554
rect 10945 -17583 24845 -17563
rect 10945 -17617 11025 -17583
rect 24765 -17617 24845 -17583
rect 10945 -17637 24845 -17617
<< mvnsubdiffcont >>
rect 11025 8733 24765 8767
rect 10965 -17557 10999 8707
rect 24791 -1906 24825 8707
rect 23145 -1979 24775 -1945
rect 23071 -6871 23105 -1995
rect 23141 -6921 24755 -6887
rect 24791 -17554 24825 -6956
rect 11025 -17617 24765 -17583
<< locali >>
rect 10965 8733 11025 8767
rect 24765 8733 24825 8767
rect 10965 8707 10999 8733
rect 24791 8707 24825 8733
rect 20173 -1651 20424 -1649
rect 19892 -1670 20424 -1651
rect 19892 -1953 20928 -1670
rect 24791 -1945 24825 -1906
rect 19892 -2094 20424 -1953
rect 23071 -1979 23145 -1945
rect 24775 -1979 24825 -1945
rect 23071 -1995 23105 -1979
rect 20164 -2345 20424 -2094
rect 20182 -2443 20424 -2345
rect 20164 -2444 20424 -2443
rect 20275 -2480 20424 -2444
rect 20275 -2548 20409 -2480
rect 17797 -3056 20814 -2895
rect 17797 -3478 18412 -3056
rect 18851 -3478 19031 -3056
rect 19470 -3478 19650 -3056
rect 20079 -3478 20259 -3056
rect 20688 -3478 20814 -3056
rect 17797 -3504 20814 -3478
rect 17797 -3505 19132 -3504
rect 17797 -3506 18491 -3505
rect 17797 -3587 17853 -3506
rect 18359 -3587 18491 -3506
rect 17797 -3732 18491 -3587
rect 18566 -3731 19132 -3505
rect 19207 -3505 20814 -3504
rect 19207 -3731 19733 -3505
rect 18566 -3732 19733 -3731
rect 19808 -3507 20814 -3505
rect 19808 -3732 20561 -3507
rect 17797 -3734 20561 -3732
rect 20636 -3734 20814 -3507
rect 17797 -3754 20814 -3734
rect 18228 -4164 18417 -3754
rect 18851 -4164 19040 -3754
rect 19456 -4164 19645 -3754
rect 20084 -4164 20273 -3754
rect 20688 -4164 20814 -3754
rect 17786 -4285 20814 -4164
rect 17689 -4549 20930 -4430
rect 18127 -4943 18263 -4549
rect 18689 -4943 18833 -4549
rect 19237 -4943 19381 -4549
rect 19807 -4943 19951 -4549
rect 20360 -4943 20504 -4549
rect 17688 -4963 20929 -4943
rect 17688 -4966 19629 -4963
rect 17688 -4967 18523 -4966
rect 17688 -5137 17952 -4967
rect 18118 -5136 18523 -4967
rect 18689 -5136 19073 -4966
rect 19239 -5133 19629 -4966
rect 19795 -5133 20187 -4963
rect 20353 -4966 20929 -4963
rect 20353 -5133 20686 -4966
rect 19239 -5136 20686 -5133
rect 20852 -5136 20929 -4966
rect 18118 -5137 20929 -5136
rect 17688 -5141 20929 -5137
rect 18132 -5544 18272 -5141
rect 18684 -5544 18828 -5141
rect 19241 -5544 19385 -5141
rect 19799 -5544 19943 -5141
rect 20356 -5544 20500 -5141
rect 17683 -5627 20932 -5544
rect 17683 -5631 19419 -5627
rect 17683 -5701 19025 -5631
rect 17683 -5805 17772 -5701
rect 18791 -5801 19025 -5701
rect 19191 -5797 19419 -5631
rect 19585 -5639 20932 -5627
rect 19585 -5797 20172 -5639
rect 19191 -5801 20172 -5797
rect 18791 -5805 20172 -5801
rect 17683 -5809 20172 -5805
rect 20338 -5809 20932 -5639
rect 17683 -5881 20932 -5809
rect 19239 -6298 19384 -5881
rect 19794 -6295 19938 -5881
rect 20360 -6295 20504 -5881
rect 24362 -2785 24809 -2683
rect 24372 -2806 24809 -2785
rect 23738 -3000 23870 -2920
rect 23738 -5906 23785 -3000
rect 23844 -5906 23870 -3000
rect 24372 -3066 24528 -2806
rect 24370 -3810 24549 -3314
rect 24451 -4505 24539 -4121
rect 24113 -4507 24886 -4505
rect 24112 -4514 24886 -4507
rect 24112 -4572 24130 -4514
rect 24683 -4572 24886 -4514
rect 24112 -4577 24886 -4572
rect 24113 -4580 24886 -4577
rect 23738 -6010 23870 -5906
rect 23546 -6260 23902 -6248
rect 23546 -6440 23728 -6260
rect 23890 -6440 23902 -6260
rect 23546 -6451 23902 -6440
rect 23071 -6887 23105 -6871
rect 23071 -6921 23141 -6887
rect 24755 -6921 24825 -6887
rect 24791 -6956 24825 -6921
rect 10965 -17583 10999 -17557
rect 24791 -17583 24825 -17554
rect 10965 -17617 11025 -17583
rect 24765 -17617 24825 -17583
<< viali >>
rect 11509 8767 24645 8788
rect 11509 8733 24645 8767
rect 11509 8722 24645 8733
rect 24770 7847 24791 8278
rect 24791 7847 24825 8278
rect 24825 7847 24845 8278
rect 10935 3390 10965 7474
rect 10965 3390 10999 7474
rect 10999 3390 11019 7474
rect 11301 3517 11336 7480
rect 20886 3498 20938 7461
rect 21189 3498 21241 7461
rect 24474 3503 24526 7466
rect 24773 3500 24791 7482
rect 24791 3500 24825 7482
rect 24825 3500 24847 7482
rect 10944 -780 10965 3184
rect 10965 -780 10999 3184
rect 10999 -780 11019 3184
rect 24771 -786 24791 3180
rect 24791 -786 24825 3180
rect 24825 -786 24845 3180
rect 10935 -6253 10965 -927
rect 10965 -6253 10999 -927
rect 10999 -6253 11022 -927
rect 24769 -1867 24791 -936
rect 24791 -1867 24825 -936
rect 24825 -1867 24844 -936
rect 23251 -1945 24717 -1928
rect 23251 -1979 24717 -1945
rect 23251 -1992 24717 -1979
rect 11385 -6348 11458 -2216
rect 19892 -2443 20182 -2345
rect 20546 -2426 20840 -2344
rect 20409 -2548 20977 -2480
rect 17853 -3587 18359 -3506
rect 18491 -3732 18566 -3505
rect 19132 -3731 19207 -3504
rect 19733 -3732 19808 -3505
rect 20561 -3734 20636 -3507
rect 17952 -5137 18118 -4967
rect 18523 -5136 18689 -4966
rect 19073 -5136 19239 -4966
rect 19629 -5133 19795 -4963
rect 20187 -5133 20353 -4963
rect 20686 -5136 20852 -4966
rect 17772 -5805 18791 -5701
rect 19025 -5801 19191 -5631
rect 19419 -5797 19585 -5627
rect 20172 -5809 20338 -5639
rect 23058 -6840 23071 -2033
rect 23071 -6840 23105 -2033
rect 23105 -6840 23118 -2033
rect 23785 -5906 23844 -3000
rect 24130 -4572 24683 -4514
rect 23728 -6440 23890 -6260
rect 23219 -6887 24656 -6868
rect 23219 -6921 24656 -6887
rect 23219 -6926 24656 -6921
rect 11246 -11938 11298 -7962
rect 24492 -11940 24544 -7964
rect 24765 -11928 24791 -7061
rect 24791 -11928 24825 -7061
rect 24825 -11928 24828 -7061
rect 10945 -16245 10965 -12264
rect 10965 -16245 10999 -12264
rect 10999 -16245 11020 -12264
rect 24772 -16242 24791 -12276
rect 24791 -16242 24825 -12276
rect 24825 -16242 24845 -12276
rect 10944 -17120 10965 -16690
rect 10965 -17120 10999 -16690
rect 10999 -17120 11019 -16690
rect 11053 -17583 24731 -17560
rect 11053 -17617 24731 -17583
rect 11053 -17636 24731 -17617
<< metal1 >>
rect 24684 8839 24905 8840
rect 11390 8788 24905 8839
rect 11390 8722 11509 8788
rect 24645 8722 24905 8788
rect 11390 8692 24905 8722
rect 10878 8624 11078 8675
rect 10878 8537 21102 8624
rect 10878 8475 11078 8537
rect 21015 8288 21102 8537
rect 11432 7856 11668 8288
rect 11764 7856 12000 8288
rect 12096 7856 12332 8288
rect 12428 7856 12664 8288
rect 12760 7856 12996 8288
rect 13092 7856 13328 8288
rect 13424 7856 13660 8288
rect 13756 7856 13992 8288
rect 14088 7856 14324 8288
rect 14420 7856 14656 8288
rect 14752 7856 14988 8288
rect 15084 7856 15320 8288
rect 15416 7856 15652 8288
rect 15748 7856 15984 8288
rect 16080 7856 16316 8288
rect 16412 7856 16648 8288
rect 16744 7856 16980 8288
rect 17076 7856 17312 8288
rect 17408 7856 17644 8288
rect 17740 7856 17976 8288
rect 18072 7856 18308 8288
rect 18404 7856 18640 8288
rect 18736 7856 18972 8288
rect 19068 7856 19304 8288
rect 19400 7856 19636 8288
rect 19732 7856 19968 8288
rect 20064 7856 20300 8288
rect 20396 7856 20632 8288
rect 20728 7856 21102 8288
rect 24684 8278 24905 8692
rect 10892 7474 11056 7509
rect 11295 7480 11342 7492
rect 10892 3390 10935 7474
rect 11019 3390 11056 7474
rect 11283 3517 11293 7480
rect 11345 3517 11355 7480
rect 20880 7461 20944 7473
rect 11295 3505 11342 3517
rect 20876 3498 20886 7461
rect 20938 3498 20948 7461
rect 20880 3486 20944 3498
rect 10892 3184 11056 3390
rect 10892 -780 10944 3184
rect 11019 -780 11056 3184
rect 10892 -927 11056 -780
rect 10892 -6253 10935 -927
rect 11022 -6253 11056 -927
rect 11432 -1779 11502 -1112
rect 11598 -1544 11834 -1112
rect 11930 -1544 12166 -1112
rect 12262 -1544 12498 -1112
rect 12594 -1544 12830 -1112
rect 12926 -1544 13162 -1112
rect 13258 -1544 13494 -1112
rect 13590 -1544 13826 -1112
rect 13922 -1544 14158 -1112
rect 14254 -1544 14490 -1112
rect 14586 -1544 14822 -1112
rect 14918 -1544 15154 -1112
rect 15250 -1544 15486 -1112
rect 15582 -1544 15818 -1112
rect 15914 -1544 16150 -1112
rect 16246 -1544 16482 -1112
rect 16578 -1544 16814 -1112
rect 16910 -1544 17146 -1112
rect 17242 -1544 17478 -1112
rect 17574 -1544 17810 -1112
rect 17906 -1544 18142 -1112
rect 18238 -1544 18474 -1112
rect 18570 -1544 18806 -1112
rect 18902 -1544 19138 -1112
rect 19234 -1544 19470 -1112
rect 19566 -1544 19802 -1112
rect 19898 -1544 20134 -1112
rect 20230 -1544 20466 -1112
rect 20562 -1544 20798 -1112
rect 11432 -1878 17362 -1779
rect 11379 -2216 11464 -2204
rect 10892 -6293 11056 -6253
rect 11375 -6348 11385 -2216
rect 11458 -6348 11468 -2216
rect 11548 -2556 11920 -2124
rect 12016 -2556 12388 -2124
rect 12484 -2556 12856 -2124
rect 12952 -2556 13324 -2124
rect 13420 -2556 13792 -2124
rect 13888 -2556 14260 -2124
rect 14356 -2556 14728 -2124
rect 14824 -2556 15196 -2124
rect 15292 -2556 15664 -2124
rect 15760 -2556 16132 -2124
rect 16228 -2556 16600 -2124
rect 16696 -2556 17068 -2124
rect 17265 -3633 17362 -1878
rect 21015 -2198 21102 7856
rect 21328 7846 21564 8278
rect 21660 7846 21896 8278
rect 21992 7846 22228 8278
rect 22324 7846 22560 8278
rect 22656 7846 22892 8278
rect 22988 7846 23224 8278
rect 23320 7846 23556 8278
rect 23652 7846 23888 8278
rect 23984 7846 24220 8278
rect 24316 7847 24770 8278
rect 24845 7847 24905 8278
rect 24316 7846 24905 7847
rect 24684 7482 24905 7846
rect 21183 7461 21247 7473
rect 24468 7466 24532 7478
rect 21179 3498 21189 7461
rect 21241 3498 21251 7461
rect 24464 3503 24474 7466
rect 24526 3503 24536 7466
rect 21183 3486 21247 3498
rect 24468 3491 24532 3503
rect 24684 3500 24773 7482
rect 24847 3500 24905 7482
rect 24684 3180 24905 3500
rect 24684 -786 24771 3180
rect 24845 -786 24905 3180
rect 24684 -936 24905 -786
rect 19985 -2266 21102 -2198
rect 21210 -1533 21382 -1468
rect 19985 -2267 21092 -2266
rect 19880 -2345 20194 -2339
rect 19880 -2443 19892 -2345
rect 20182 -2443 20194 -2345
rect 20534 -2344 20852 -2338
rect 20534 -2426 20546 -2344
rect 20840 -2426 20852 -2344
rect 20534 -2432 20852 -2426
rect 19880 -2449 20194 -2443
rect 19901 -2658 20162 -2449
rect 20397 -2480 20989 -2474
rect 20397 -2548 20409 -2480
rect 20977 -2548 20989 -2480
rect 20397 -2554 20989 -2548
rect 20488 -2658 20862 -2554
rect 19901 -2875 20855 -2658
rect 19901 -2876 20162 -2875
rect 20845 -2876 20855 -2875
rect 20923 -2876 20933 -2658
rect 20881 -3060 20949 -3050
rect 19870 -3172 20294 -3171
rect 18584 -3223 20294 -3172
rect 20440 -3218 20881 -3176
rect 18584 -3224 19920 -3223
rect 18507 -3489 18553 -3276
rect 17841 -3506 18371 -3500
rect 17841 -3587 17853 -3506
rect 18359 -3587 18371 -3506
rect 17841 -3593 18371 -3587
rect 18344 -3633 18388 -3631
rect 17265 -3677 18388 -3633
rect 17265 -5541 17362 -3677
rect 17799 -3946 17954 -3902
rect 17799 -4088 17843 -3946
rect 17908 -4053 18071 -4012
rect 17770 -4272 17780 -4088
rect 17845 -4272 17855 -4088
rect 17789 -4278 17843 -4272
rect 17524 -4536 17534 -4378
rect 17593 -4536 17603 -4378
rect 17540 -5418 17589 -4536
rect 17789 -4828 17832 -4278
rect 17908 -4286 17949 -4053
rect 17899 -4444 17909 -4286
rect 17968 -4444 17978 -4286
rect 18107 -4440 18182 -3879
rect 18344 -3901 18388 -3677
rect 18449 -3725 18459 -3489
rect 18622 -3725 18632 -3489
rect 18485 -3732 18491 -3725
rect 18566 -3732 18572 -3725
rect 18485 -3744 18572 -3732
rect 18344 -3945 18564 -3901
rect 17908 -4450 17949 -4444
rect 18061 -4601 18071 -4440
rect 18228 -4601 18238 -4440
rect 17877 -4681 18218 -4659
rect 17877 -4700 18169 -4681
rect 18007 -4858 18057 -4739
rect 18159 -4848 18169 -4700
rect 18226 -4848 18236 -4681
rect 18344 -4820 18388 -3945
rect 18728 -3968 18769 -3280
rect 19148 -3492 19194 -3277
rect 19126 -3494 19213 -3492
rect 19080 -3730 19090 -3494
rect 19253 -3730 19263 -3494
rect 19126 -3731 19132 -3730
rect 19207 -3731 19213 -3730
rect 19126 -3743 19213 -3731
rect 18612 -4188 18653 -4021
rect 19125 -4188 19169 -3878
rect 19354 -3968 19395 -3280
rect 19745 -3493 19791 -3279
rect 19727 -3502 19814 -3493
rect 19683 -3738 19693 -3502
rect 19856 -3738 19866 -3502
rect 19727 -3744 19814 -3738
rect 18612 -4232 19169 -4188
rect 19236 -4193 19277 -4019
rect 19725 -4193 19769 -3879
rect 19953 -3965 19994 -3277
rect 20242 -3296 20294 -3223
rect 20881 -3247 20949 -3237
rect 20242 -3344 20425 -3296
rect 20242 -3903 20294 -3344
rect 20577 -3495 20626 -3280
rect 21021 -3333 21075 -2267
rect 21210 -2350 21275 -1533
rect 21494 -1554 21730 -1122
rect 21826 -1554 22062 -1122
rect 22158 -1554 22394 -1122
rect 22490 -1554 22726 -1122
rect 22822 -1554 23058 -1122
rect 23154 -1554 23390 -1122
rect 23486 -1554 23722 -1122
rect 23818 -1554 24054 -1122
rect 24150 -1554 24386 -1122
rect 24684 -1812 24769 -936
rect 22994 -1867 24769 -1812
rect 24844 -1867 24905 -936
rect 22994 -1928 24905 -1867
rect 22994 -1992 23251 -1928
rect 24717 -1992 24905 -1928
rect 22994 -2033 24905 -1992
rect 21414 -2212 21424 -2054
rect 22870 -2212 22880 -2054
rect 20829 -3387 21075 -3333
rect 21150 -2466 21275 -2350
rect 20555 -3500 20642 -3495
rect 20507 -3736 20517 -3500
rect 20680 -3736 20690 -3500
rect 20555 -3746 20642 -3736
rect 20242 -3947 20418 -3903
rect 20242 -3952 20406 -3947
rect 18612 -4280 18653 -4232
rect 18457 -4338 18467 -4280
rect 18653 -4338 18663 -4280
rect 18465 -4692 18506 -4338
rect 18562 -4858 18612 -4738
rect 18915 -4818 18959 -4232
rect 19236 -4237 19769 -4193
rect 19236 -4288 19277 -4237
rect 19017 -4329 19277 -4288
rect 19017 -4689 19058 -4329
rect 17787 -4908 18057 -4858
rect 18337 -4908 18612 -4858
rect 19111 -4861 19161 -4737
rect 19469 -4828 19513 -4237
rect 19848 -4312 19889 -4021
rect 20242 -4025 20294 -3952
rect 20577 -3973 20626 -3746
rect 20242 -4077 20535 -4025
rect 19848 -4323 19925 -4312
rect 19580 -4364 19925 -4323
rect 19580 -4689 19621 -4364
rect 19851 -4375 19925 -4364
rect 20148 -4375 20158 -4312
rect 19670 -4861 19720 -4741
rect 17787 -5365 17837 -4908
rect 17946 -4967 18124 -4955
rect 17946 -5137 17952 -4967
rect 18118 -5137 18124 -4967
rect 17946 -5149 18124 -5137
rect 18009 -5360 18061 -5149
rect 18337 -5365 18387 -4908
rect 18897 -4911 19161 -4861
rect 19461 -4911 19720 -4861
rect 18517 -4966 18695 -4954
rect 18517 -5136 18523 -4966
rect 18689 -5136 18695 -4966
rect 18517 -5148 18695 -5136
rect 18573 -5362 18625 -5148
rect 18897 -5364 18947 -4911
rect 19067 -4966 19245 -4954
rect 19067 -5136 19073 -4966
rect 19239 -5136 19245 -4966
rect 19067 -5148 19245 -5136
rect 19127 -5364 19179 -5148
rect 19461 -5364 19511 -4911
rect 19623 -4963 19801 -4951
rect 19623 -5133 19629 -4963
rect 19795 -5133 19801 -4963
rect 19623 -5145 19801 -5133
rect 19681 -5366 19733 -5145
rect 19851 -5169 19892 -4375
rect 20242 -4498 20294 -4077
rect 20383 -4377 20393 -4314
rect 20616 -4319 20626 -4314
rect 20829 -4319 20883 -3387
rect 21150 -3618 21215 -2466
rect 21257 -3266 21267 -3089
rect 21335 -3206 21345 -3089
rect 21646 -3150 22088 -3089
rect 21646 -3206 21707 -3150
rect 21335 -3266 21707 -3206
rect 21274 -3267 21707 -3266
rect 21080 -3689 21215 -3618
rect 21277 -3606 21426 -3544
rect 20932 -4108 20942 -3836
rect 21017 -4108 21027 -3836
rect 20616 -4373 20883 -4319
rect 20616 -4377 20626 -4373
rect 20001 -4550 20294 -4498
rect 20001 -4816 20053 -4550
rect 20951 -4643 21005 -4108
rect 20102 -4673 21005 -4643
rect 20102 -4697 20400 -4673
rect 20217 -4861 20267 -4745
rect 20390 -4840 20400 -4697
rect 20457 -4697 21005 -4673
rect 20457 -4840 20467 -4697
rect 20005 -4911 20267 -4861
rect 19830 -5346 19840 -5169
rect 19911 -5346 19921 -5169
rect 20005 -5366 20055 -4911
rect 20181 -4963 20359 -4951
rect 20181 -5133 20187 -4963
rect 20353 -5133 20359 -4963
rect 20181 -5145 20359 -5133
rect 20242 -5357 20294 -5145
rect 17540 -5467 17964 -5418
rect 20562 -5421 20619 -4739
rect 21080 -4749 21145 -3689
rect 20767 -4811 21005 -4751
rect 20680 -4966 20858 -4954
rect 20680 -5136 20686 -4966
rect 20852 -5136 20858 -4966
rect 20680 -5148 20858 -5136
rect 20791 -5364 20851 -5148
rect 18432 -5479 20735 -5421
rect 17265 -5580 18950 -5541
rect 11379 -6360 11464 -6348
rect 10878 -6538 11078 -6495
rect 10878 -6645 11564 -6538
rect 10878 -6695 11078 -6645
rect 11782 -6756 12154 -6324
rect 12250 -6756 12622 -6324
rect 12718 -6756 13090 -6324
rect 13186 -6756 13558 -6324
rect 13654 -6756 14026 -6324
rect 14122 -6756 14494 -6324
rect 14590 -6756 14962 -6324
rect 15058 -6756 15430 -6324
rect 15526 -6756 15898 -6324
rect 15994 -6756 16366 -6324
rect 16462 -6756 16834 -6324
rect 17265 -6490 17362 -5580
rect 17760 -5701 18803 -5695
rect 17760 -5805 17772 -5701
rect 18791 -5805 18803 -5701
rect 17760 -5811 18803 -5805
rect 18911 -6091 18950 -5580
rect 19019 -5631 19197 -5619
rect 19413 -5627 19591 -5615
rect 19015 -5801 19025 -5631
rect 19191 -5801 19201 -5631
rect 19409 -5797 19419 -5627
rect 19585 -5797 19595 -5627
rect 19831 -5797 19841 -5620
rect 19912 -5797 19922 -5620
rect 19019 -5813 19197 -5801
rect 19413 -5809 19591 -5797
rect 19126 -6093 19178 -5813
rect 19459 -6091 19511 -5809
rect 19842 -6016 19890 -5797
rect 19670 -6064 19890 -6016
rect 20022 -6083 20066 -5479
rect 20166 -5639 20344 -5627
rect 20162 -5809 20172 -5639
rect 20338 -5809 20348 -5639
rect 20166 -5821 20344 -5809
rect 20224 -6089 20276 -5821
rect 20580 -6079 20635 -5479
rect 20670 -5775 20678 -5707
rect 20878 -5775 20888 -5707
rect 20787 -6084 20837 -5775
rect 18984 -6143 20550 -6136
rect 18984 -6192 20485 -6143
rect 20475 -6320 20485 -6192
rect 20556 -6320 20566 -6143
rect 20494 -6327 20550 -6320
rect 20680 -6367 20732 -6134
rect 20670 -6435 20680 -6367
rect 20880 -6435 20890 -6367
rect 17049 -6612 17362 -6490
rect 20945 -7032 21005 -4811
rect 21060 -4803 21145 -4749
rect 21060 -5700 21125 -4803
rect 21277 -4855 21339 -3606
rect 21385 -4045 21579 -4040
rect 21381 -4243 21391 -4045
rect 21573 -4243 21583 -4045
rect 22994 -4118 23058 -2033
rect 21173 -4915 21339 -4855
rect 21385 -4668 21579 -4243
rect 21385 -4860 21396 -4668
rect 21575 -4860 21585 -4668
rect 22846 -4794 23058 -4118
rect 21385 -4869 21579 -4860
rect 21045 -5712 21136 -5700
rect 21045 -5889 21055 -5712
rect 21126 -5889 21136 -5712
rect 21173 -5983 21233 -4915
rect 21073 -6043 21233 -5983
rect 21282 -5126 21437 -5066
rect 21073 -6099 21133 -6043
rect 21055 -6276 21065 -6099
rect 21136 -6276 21146 -6099
rect 21282 -6370 21342 -5126
rect 21100 -6438 21110 -6370
rect 21310 -6437 21342 -6370
rect 21310 -6438 21320 -6437
rect 21422 -6871 21432 -6710
rect 22858 -6871 22868 -6710
rect 22994 -6840 23058 -4794
rect 23118 -6793 23219 -2033
rect 24712 -2262 24912 -2207
rect 23525 -2339 24912 -2262
rect 23525 -3162 23602 -2339
rect 24712 -2407 24912 -2339
rect 23716 -2586 24446 -2568
rect 23716 -2756 24260 -2586
rect 24425 -2756 24446 -2586
rect 23716 -2770 24446 -2756
rect 23716 -3000 23936 -2770
rect 23329 -5840 23339 -5786
rect 23454 -5840 23464 -5786
rect 23402 -6414 23454 -5840
rect 23514 -6554 23612 -5852
rect 23716 -5906 23785 -3000
rect 23844 -4297 23936 -3000
rect 24474 -2952 24698 -2903
rect 24474 -3181 24523 -2952
rect 24458 -3238 24468 -3181
rect 24527 -3238 24538 -3181
rect 24590 -3774 24643 -3430
rect 24472 -3974 24643 -3774
rect 24683 -4035 24723 -3701
rect 24266 -4075 24723 -4035
rect 23966 -4266 23976 -4214
rect 24066 -4215 24076 -4214
rect 24266 -4215 24308 -4075
rect 24066 -4225 24308 -4215
rect 24066 -4255 24270 -4225
rect 24066 -4266 24076 -4255
rect 24468 -4257 24478 -4205
rect 24530 -4217 24540 -4205
rect 24530 -4257 24727 -4217
rect 23844 -4389 24255 -4297
rect 24342 -4358 24667 -4313
rect 23844 -4506 24024 -4389
rect 23844 -4514 24696 -4506
rect 23844 -4572 24130 -4514
rect 24683 -4572 24696 -4514
rect 23844 -4582 24696 -4572
rect 23844 -4753 24024 -4582
rect 24343 -4725 24353 -4670
rect 24407 -4680 24417 -4670
rect 24407 -4714 24725 -4680
rect 24407 -4725 24417 -4714
rect 23844 -4840 24678 -4753
rect 23844 -5906 23936 -4840
rect 24760 -4876 24859 -3423
rect 24545 -4974 24859 -4876
rect 23716 -6219 23936 -5906
rect 23716 -6260 24444 -6219
rect 23716 -6440 23728 -6260
rect 23890 -6440 24444 -6260
rect 23716 -6451 24444 -6440
rect 24545 -6554 24643 -4974
rect 23514 -6652 24643 -6554
rect 23118 -6840 24882 -6793
rect 22994 -6868 24882 -6840
rect 22994 -6926 23219 -6868
rect 24656 -6926 24882 -6868
rect 22994 -6934 24882 -6926
rect 22995 -6944 24882 -6934
rect 20945 -7092 24406 -7032
rect 11388 -7722 11625 -7290
rect 11719 -7722 11956 -7290
rect 12050 -7722 12287 -7290
rect 12381 -7722 12618 -7290
rect 12712 -7722 12949 -7290
rect 13043 -7722 13280 -7290
rect 13374 -7722 13611 -7290
rect 13705 -7722 13942 -7290
rect 14036 -7722 14273 -7290
rect 14367 -7722 14604 -7290
rect 14698 -7722 14935 -7290
rect 15029 -7722 15266 -7290
rect 15360 -7722 15597 -7290
rect 15691 -7722 15928 -7290
rect 16022 -7722 16259 -7290
rect 16353 -7722 16590 -7290
rect 16684 -7722 16921 -7290
rect 17015 -7722 17252 -7290
rect 17346 -7722 17583 -7290
rect 17677 -7722 17914 -7290
rect 18008 -7722 18245 -7290
rect 18339 -7722 18576 -7290
rect 18670 -7722 18907 -7290
rect 19001 -7722 19238 -7290
rect 19332 -7722 19569 -7290
rect 19663 -7722 19900 -7290
rect 19994 -7722 20231 -7290
rect 20325 -7722 20562 -7290
rect 20656 -7722 20893 -7290
rect 20987 -7722 21224 -7290
rect 21318 -7722 21555 -7290
rect 21649 -7722 21886 -7290
rect 21980 -7722 22217 -7290
rect 22311 -7722 22548 -7290
rect 22642 -7722 22879 -7290
rect 22973 -7722 23210 -7290
rect 23304 -7722 23541 -7290
rect 23635 -7722 23872 -7290
rect 23966 -7722 24203 -7290
rect 24336 -7722 24406 -7092
rect 24731 -7061 24882 -6944
rect 11240 -7962 11304 -7950
rect 11236 -11938 11246 -7962
rect 11298 -11938 11308 -7962
rect 24486 -7964 24550 -7952
rect 11240 -11950 11304 -11938
rect 24482 -11940 24492 -7964
rect 24544 -11940 24554 -7964
rect 24731 -11928 24765 -7061
rect 24828 -11928 24882 -7061
rect 24486 -11952 24550 -11940
rect 10939 -12264 11026 -12252
rect 10935 -16245 10945 -12264
rect 11020 -16245 11030 -12264
rect 24731 -12276 24882 -11928
rect 24731 -16242 24772 -12276
rect 24845 -16242 24882 -12276
rect 10938 -16257 11026 -16245
rect 10938 -16690 11025 -16257
rect 10938 -17120 10944 -16690
rect 11019 -17120 11458 -16690
rect 10938 -17122 11458 -17120
rect 11554 -17122 11790 -16690
rect 11886 -17122 12122 -16690
rect 12218 -17122 12454 -16690
rect 12550 -17122 12786 -16690
rect 12882 -17122 13118 -16690
rect 13214 -17122 13450 -16690
rect 13546 -17122 13782 -16690
rect 13878 -17122 14114 -16690
rect 14210 -17122 14446 -16690
rect 14542 -17122 14778 -16690
rect 14874 -17122 15110 -16690
rect 15206 -17122 15442 -16690
rect 15538 -17122 15774 -16690
rect 15870 -17122 16106 -16690
rect 16202 -17122 16438 -16690
rect 16534 -17122 16770 -16690
rect 16866 -17122 17102 -16690
rect 17198 -17122 17434 -16690
rect 17530 -17122 17766 -16690
rect 17862 -17122 18098 -16690
rect 18194 -17122 18430 -16690
rect 18526 -17122 18762 -16690
rect 18858 -17122 19094 -16690
rect 19190 -17122 19426 -16690
rect 19522 -17122 19758 -16690
rect 19854 -17122 20090 -16690
rect 20186 -17122 20422 -16690
rect 20518 -17122 20754 -16690
rect 20850 -17122 21086 -16690
rect 21182 -17122 21418 -16690
rect 21514 -17122 21750 -16690
rect 21846 -17122 22082 -16690
rect 22178 -17122 22414 -16690
rect 22510 -17122 22746 -16690
rect 22842 -17122 23078 -16690
rect 23174 -17122 23410 -16690
rect 23506 -17122 23742 -16690
rect 23838 -17122 24074 -16690
rect 24170 -17122 24406 -16690
rect 10938 -17132 11025 -17122
rect 24731 -17485 24882 -16242
rect 10903 -17560 24882 -17485
rect 10903 -17636 11053 -17560
rect 24731 -17636 24882 -17560
rect 10903 -17688 24882 -17636
<< via1 >>
rect 11293 3517 11301 7480
rect 11301 3517 11336 7480
rect 11336 3517 11345 7480
rect 20886 3498 20938 7461
rect 10944 -780 11019 3184
rect 11385 -6348 11458 -2216
rect 21189 3498 21241 7461
rect 24474 3503 24526 7466
rect 24771 -786 24845 3180
rect 20546 -2426 20792 -2344
rect 20855 -2876 20923 -2658
rect 17853 -3587 18359 -3506
rect 17780 -4272 17845 -4088
rect 17534 -4536 17593 -4378
rect 17909 -4444 17968 -4286
rect 18459 -3505 18622 -3489
rect 18459 -3725 18491 -3505
rect 18491 -3725 18566 -3505
rect 18566 -3725 18622 -3505
rect 18071 -4601 18228 -4440
rect 18169 -4848 18226 -4681
rect 19090 -3504 19253 -3494
rect 19090 -3730 19132 -3504
rect 19132 -3730 19207 -3504
rect 19207 -3730 19253 -3504
rect 19693 -3505 19856 -3502
rect 19693 -3732 19733 -3505
rect 19733 -3732 19808 -3505
rect 19808 -3732 19856 -3505
rect 19693 -3738 19856 -3732
rect 20881 -3237 20949 -3060
rect 21424 -2212 22870 -2054
rect 20517 -3507 20680 -3500
rect 20517 -3734 20561 -3507
rect 20561 -3734 20636 -3507
rect 20636 -3734 20680 -3507
rect 20517 -3736 20680 -3734
rect 18467 -4338 18653 -4280
rect 19925 -4375 20148 -4312
rect 20393 -4377 20616 -4314
rect 21267 -3266 21335 -3089
rect 20942 -4108 21017 -3836
rect 20400 -4840 20457 -4673
rect 19840 -5346 19911 -5169
rect 17772 -5805 18791 -5701
rect 19025 -5801 19191 -5631
rect 19419 -5797 19585 -5627
rect 19841 -5797 19912 -5620
rect 20172 -5809 20338 -5639
rect 20678 -5775 20878 -5707
rect 20485 -6320 20556 -6143
rect 20680 -6435 20880 -6367
rect 21391 -4243 21573 -4045
rect 21396 -4860 21575 -4668
rect 21055 -5889 21126 -5712
rect 21065 -6276 21136 -6099
rect 21110 -6438 21310 -6370
rect 21432 -6871 22858 -6710
rect 24260 -2756 24425 -2586
rect 23339 -5840 23454 -5786
rect 24468 -3238 24527 -3181
rect 24018 -3952 24253 -3794
rect 23976 -4266 24066 -4214
rect 24478 -4257 24530 -4205
rect 24353 -4725 24407 -4670
rect 24290 -5129 24455 -4959
rect 11246 -11938 11298 -7962
rect 24492 -11940 24544 -7964
rect 10945 -16245 11020 -12264
rect 24772 -16242 24845 -12276
<< metal2 >>
rect 11293 7489 11345 7490
rect 10878 7480 24912 7489
rect 10878 3517 11293 7480
rect 11345 7466 24912 7480
rect 11345 7461 24474 7466
rect 11345 3517 20886 7461
rect 10878 3498 20886 3517
rect 20938 3498 21189 7461
rect 21241 3503 24474 7461
rect 24526 3503 24912 7466
rect 21241 3498 24912 3503
rect 10878 3489 24912 3498
rect 20886 3488 20938 3489
rect 21189 3488 21241 3489
rect 10878 3184 24912 3204
rect 10878 -780 10944 3184
rect 11019 3180 24912 3184
rect 11019 -780 24771 3180
rect 10878 -786 24771 -780
rect 24845 -786 24912 3180
rect 10878 -796 24912 -786
rect 11301 -2216 11505 -2088
rect 11301 -6348 11385 -2216
rect 11458 -2677 11505 -2216
rect 11458 -6189 17081 -2677
rect 17536 -3380 18742 -796
rect 19713 -1989 20919 -796
rect 19713 -2344 20792 -1989
rect 19713 -2426 20546 -2344
rect 19713 -3380 20792 -2426
rect 21392 -2054 22883 -1618
rect 21392 -2212 21424 -2054
rect 22870 -2212 22883 -2054
rect 21392 -2224 22883 -2212
rect 20855 -2658 20923 -2648
rect 21392 -2658 21588 -2224
rect 20923 -2875 21588 -2658
rect 23980 -2586 24912 -2570
rect 23980 -2756 24260 -2586
rect 24425 -2756 24912 -2586
rect 23980 -2770 24912 -2756
rect 20855 -2886 20923 -2876
rect 20871 -3237 20881 -3060
rect 20949 -3157 20959 -3060
rect 21267 -3089 21335 -3079
rect 20949 -3237 21267 -3157
rect 20871 -3244 21267 -3237
rect 20871 -3247 21016 -3244
rect 17536 -3489 20792 -3380
rect 17536 -3506 18459 -3489
rect 17536 -3587 17853 -3506
rect 18359 -3587 18459 -3506
rect 17536 -3725 18459 -3587
rect 18622 -3494 20792 -3489
rect 18622 -3725 19090 -3494
rect 17536 -3730 19090 -3725
rect 19253 -3500 20792 -3494
rect 19253 -3502 20517 -3500
rect 19253 -3730 19693 -3502
rect 17536 -3738 19693 -3730
rect 19856 -3736 20517 -3502
rect 20680 -3736 20792 -3500
rect 19856 -3738 20792 -3736
rect 17536 -3827 20792 -3738
rect 20942 -3830 21016 -3247
rect 21267 -3276 21335 -3266
rect 20942 -3836 21017 -3830
rect 17780 -4088 17845 -4078
rect 21392 -4035 21588 -2875
rect 23898 -3000 24407 -2946
rect 23992 -3778 24273 -3776
rect 23992 -3794 24289 -3778
rect 23992 -3952 24018 -3794
rect 24253 -3952 24289 -3794
rect 23992 -3974 24289 -3952
rect 20942 -4118 21017 -4108
rect 21391 -4045 21588 -4035
rect 17845 -4205 20734 -4153
rect 17780 -4282 17845 -4272
rect 17909 -4286 17968 -4276
rect 17534 -4378 17593 -4368
rect 17593 -4427 17909 -4382
rect 18467 -4280 18653 -4270
rect 17968 -4333 18467 -4288
rect 20682 -4295 20734 -4205
rect 21573 -4243 21588 -4045
rect 23976 -4214 24066 -4204
rect 21391 -4244 21588 -4243
rect 21391 -4253 21573 -4244
rect 23267 -4266 23976 -4215
rect 23267 -4267 24066 -4266
rect 23267 -4295 23319 -4267
rect 23976 -4275 24066 -4267
rect 18467 -4348 18653 -4338
rect 19925 -4306 20148 -4302
rect 20393 -4306 20616 -4304
rect 19925 -4312 20616 -4306
rect 20148 -4314 20616 -4312
rect 20148 -4375 20393 -4314
rect 19925 -4377 20393 -4375
rect 20682 -4347 23319 -4295
rect 19925 -4381 20616 -4377
rect 19925 -4385 20148 -4381
rect 20393 -4387 20616 -4381
rect 18071 -4440 18228 -4430
rect 24123 -4440 24289 -3974
rect 17909 -4454 17968 -4444
rect 17534 -4546 17593 -4536
rect 18062 -4601 18071 -4440
rect 18228 -4601 24289 -4440
rect 18071 -4611 18228 -4601
rect 18169 -4681 18226 -4671
rect 20400 -4673 20457 -4663
rect 18226 -4751 20400 -4690
rect 18169 -4858 18226 -4848
rect 20400 -4850 20457 -4840
rect 21396 -4667 21575 -4658
rect 21396 -4668 21580 -4667
rect 21575 -4860 21580 -4668
rect 21396 -4870 21580 -4860
rect 19840 -5169 19911 -5159
rect 19840 -5356 19911 -5346
rect 17535 -5627 19646 -5594
rect 19849 -5610 19897 -5356
rect 17535 -5631 19419 -5627
rect 17535 -5701 19025 -5631
rect 17535 -5805 17772 -5701
rect 18791 -5801 19025 -5701
rect 19191 -5797 19419 -5631
rect 19585 -5797 19646 -5627
rect 19191 -5801 19646 -5797
rect 18791 -5805 19646 -5801
rect 17535 -6067 19646 -5805
rect 19841 -5620 19912 -5610
rect 19841 -5807 19912 -5797
rect 19991 -5639 20387 -5597
rect 19991 -5809 20172 -5639
rect 20338 -5809 20387 -5639
rect 20678 -5702 20878 -5697
rect 21055 -5702 21126 -5700
rect 20678 -5707 21126 -5702
rect 20878 -5712 21126 -5707
rect 20878 -5775 21055 -5712
rect 20678 -5785 20878 -5775
rect 19991 -6067 20387 -5809
rect 21055 -5900 21126 -5889
rect 11458 -6348 11505 -6189
rect 11301 -7948 11505 -6348
rect 17535 -6620 20387 -6067
rect 21065 -6099 21136 -6089
rect 20485 -6143 20556 -6133
rect 20556 -6232 21065 -6170
rect 21065 -6286 21136 -6276
rect 20485 -6330 20556 -6320
rect 20680 -6367 20880 -6357
rect 21110 -6370 21310 -6360
rect 20880 -6432 21110 -6374
rect 20680 -6445 20880 -6435
rect 21110 -6448 21310 -6438
rect 17535 -7948 18741 -6620
rect 19708 -6753 20387 -6620
rect 21403 -6673 21580 -4870
rect 24123 -4945 24289 -4601
rect 24353 -4670 24407 -3000
rect 24468 -3181 24527 -3171
rect 24712 -3181 24912 -3047
rect 24527 -3238 24912 -3181
rect 24468 -3248 24527 -3238
rect 24712 -3247 24912 -3238
rect 24478 -4195 24517 -3248
rect 24478 -4205 24530 -4195
rect 24478 -4267 24530 -4257
rect 24478 -4275 24517 -4267
rect 24353 -4738 24407 -4725
rect 24123 -4959 24455 -4945
rect 24123 -5129 24290 -4959
rect 24455 -5129 24912 -5045
rect 24123 -5245 24912 -5129
rect 24712 -5599 24912 -5530
rect 24125 -5653 24912 -5599
rect 24712 -5730 24912 -5653
rect 23339 -5786 23454 -5776
rect 23339 -5850 23454 -5840
rect 21403 -6710 22888 -6673
rect 19708 -7948 20914 -6753
rect 21403 -6871 21432 -6710
rect 22858 -6871 22888 -6710
rect 21403 -7948 22888 -6871
rect 10878 -7962 24912 -7948
rect 10878 -11938 11246 -7962
rect 11298 -7964 24912 -7962
rect 11298 -11938 24492 -7964
rect 10878 -11940 24492 -11938
rect 24544 -11940 24912 -7964
rect 10878 -11948 24912 -11940
rect 24492 -11950 24544 -11948
rect 10945 -12256 11020 -12254
rect 10878 -12264 24912 -12256
rect 10878 -16245 10945 -12264
rect 11020 -12276 24912 -12264
rect 11020 -16242 24772 -12276
rect 24845 -16242 24912 -12276
rect 11020 -16245 24912 -16242
rect 10878 -16256 24912 -16245
use sky130_fd_pr__diode_pd2nw_05v5_K4SERG  D1
timestamp 1698702074
transform 1 0 20692 0 1 -2231
box -321 -321 321 321
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D2
timestamp 1698702074
transform 1 0 20038 0 1 -2234
box -183 -183 183 183
use level_shifter  level_shifter_0
timestamp 1698861938
transform -1 0 24050 0 -1 -4485
box -422 -2464 2736 144
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  sky130_fd_pr__diode_pw2nd_05v5_FT76RJ_0
timestamp 1698702074
transform 1 0 24663 0 1 -2920
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  sky130_fd_pr__diode_pw2nd_05v5_FT76RJ_1
timestamp 1698702074
transform 1 0 23433 0 1 -6395
box -183 -183 183 183
use sky130_fd_pr__pfet_01v8_LGS3BL  sky130_fd_pr__pfet_01v8_LGS3BL_0
timestamp 1698716925
transform -1 0 24701 0 1 -3562
box -211 -284 211 284
use level_shifter  x2
timestamp 1698861938
transform -1 0 24050 0 1 -4413
box -422 -2464 2736 144
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM1
timestamp 1698788623
transform -1 0 19592 0 1 -4751
box -278 -269 278 269
use sky130_fd_pr__pfet_g5v0d10v5_XHZHTH  XM2
timestamp 1698788623
transform -1 0 19868 0 1 -3960
box -308 -304 308 304
use sky130_fd_pr__pfet_g5v0d10v5_XHZHTH  XM3
timestamp 1698788623
transform -1 0 19252 0 1 -3960
box -308 -304 308 304
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM4
timestamp 1698788623
transform -1 0 19036 0 1 -4751
box -278 -269 278 269
use sky130_fd_pr__nfet_01v8_L9WNCD  XM5
timestamp 1698716925
transform -1 0 24288 0 -1 -4313
box -211 -229 211 229
use sky130_fd_pr__pfet_g5v0d10v5_XHZHTH  XM9
timestamp 1698788623
transform -1 0 18636 0 1 -3960
box -308 -304 308 304
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM10
timestamp 1698788623
transform -1 0 18480 0 1 -4751
box -278 -269 278 269
use sky130_fd_pr__pfet_g5v0d10v5_XHZHTH  XM11
timestamp 1698788623
transform -1 0 18020 0 1 -3960
box -308 -304 308 304
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM12
timestamp 1698788623
transform -1 0 17924 0 -1 -5351
box -278 -269 278 269
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM13
timestamp 1698788623
transform -1 0 17924 0 1 -4751
box -278 -269 278 269
use sky130_fd_pr__nfet_01v8_L9KS9E  XM14
timestamp 1698716925
transform -1 0 24701 0 1 -4313
box -211 -229 211 229
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM21
timestamp 1698788623
transform -1 0 20704 0 -1 -5351
box -278 -269 278 269
use sky130_fd_pr__pfet_g5v0d10v5_XHZHTH  XM22
timestamp 1698788623
transform -1 0 20484 0 1 -3960
box -308 -304 308 304
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM23
timestamp 1698788623
transform -1 0 20704 0 1 -4751
box -278 -269 278 269
use sky130_fd_pr__pfet_g5v0d10v5_XHZHTH  XM24
timestamp 1698788623
transform -1 0 19868 0 -1 -3282
box -308 -304 308 304
use sky130_fd_pr__pfet_g5v0d10v5_XHZHTH  XM25
timestamp 1698788623
transform -1 0 19252 0 -1 -3282
box -308 -304 308 304
use sky130_fd_pr__pfet_g5v0d10v5_XHZHTH  XM26
timestamp 1698788623
transform -1 0 18636 0 -1 -3282
box -308 -304 308 304
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM27
timestamp 1698788623
transform -1 0 18480 0 -1 -5351
box -278 -269 278 269
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM28
timestamp 1698788623
transform -1 0 19036 0 -1 -5351
box -278 -269 278 269
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM29
timestamp 1698788623
transform -1 0 19592 0 -1 -5351
box -278 -269 278 269
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM30
timestamp 1698788623
transform -1 0 20148 0 -1 -5351
box -278 -269 278 269
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM31
timestamp 1698788623
transform -1 0 19594 0 -1 -6077
box -278 -269 278 269
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM32
timestamp 1698788623
transform -1 0 19038 0 -1 -6077
box -278 -269 278 269
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM33
timestamp 1698788623
transform -1 0 20150 0 -1 -6077
box -278 -269 278 269
use sky130_fd_pr__pfet_g5v0d10v5_XHZHTH  XM34
timestamp 1698788623
transform -1 0 20484 0 -1 -3282
box -308 -304 308 304
use sky130_fd_pr__nfet_01v8_L78EGD  XM35
timestamp 1698716925
transform -1 0 24701 0 1 -4763
box -211 -221 211 221
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM36
timestamp 1698788623
transform -1 0 20148 0 1 -4751
box -278 -269 278 269
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM46
timestamp 1698788623
transform -1 0 20706 0 -1 -6077
box -278 -269 278 269
use sky130_fd_pr__res_xhigh_po_0p35_6T4SHR  XR1
timestamp 1698702074
transform 1 0 17897 0 1 -12206
box -6675 -5082 6675 5082
use sky130_fd_pr__res_high_po_0p69_7CN4E3  XR2
timestamp 1698702074
transform 1 0 14308 0 1 -4440
box -2926 -2482 2926 2482
use sky130_fd_pr__res_xhigh_po_0p35_6T4E5R  XR3
timestamp 1698702074
transform -1 0 16115 0 1 3372
box -4849 -5082 4849 5082
use sky130_fd_pr__res_xhigh_po_0p35_9AHPBN  XR4
timestamp 1698702074
transform -1 0 22857 0 1 3362
box -1695 -5082 1695 5082
use sky130_fd_pr__res_high_po_0p69_CY6CB8  XR8
timestamp 1698702074
transform -1 0 23565 0 -1 -4466
box -235 -1582 235 1582
<< labels >>
flabel metal1 10878 -6695 11078 -6495 0 FreeSans 800 0 0 0 out
port 1 nsew
flabel metal1 10878 8475 11078 8675 0 FreeSans 800 0 0 0 in
port 0 nsew
flabel metal1 24712 -2407 24912 -2207 0 FreeSans 800 0 0 0 dout
port 7 nsew
flabel metal2 24712 -2770 24912 -2570 0 FreeSans 800 0 0 0 dvss
port 4 nsew
flabel metal2 24712 -3247 24912 -3047 0 FreeSans 800 0 0 0 ena
port 6 nsew
flabel metal2 24712 -5245 24912 -5045 0 FreeSans 800 0 0 0 dvdd
port 5 nsew
flabel metal2 24712 -5730 24912 -5530 0 FreeSans 800 0 0 0 boost
port 8 nsew
flabel metal2 s 10878 -796 11220 3204 0 FreeSans 1280 90 0 0 avdd
port 2 nsew
flabel metal2 10878 -11948 11220 -7948 0 FreeSans 1280 90 0 0 avss
port 3 nsew
flabel metal2 24570 -11948 24912 -7948 0 FreeSans 1280 90 0 0 avss
port 3 nsew
flabel metal2 10878 3489 11220 7489 0 FreeSans 1280 90 0 0 avss
port 3 nsew
flabel metal2 24570 3489 24912 7489 0 FreeSans 1280 90 0 0 avss
port 3 nsew
flabel metal2 s 24570 -796 24912 3204 0 FreeSans 1280 90 0 0 avdd
port 2 nsew
flabel metal2 s 10878 -16256 11220 -12256 0 FreeSans 1280 90 0 0 avdd
port 2 nsew
flabel metal2 s 24570 -16256 24912 -12256 0 FreeSans 1280 90 0 0 avdd
port 2 nsew
<< end >>
