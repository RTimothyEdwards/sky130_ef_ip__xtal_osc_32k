magic
tech sky130A
magscale 1 2
timestamp 1698702074
<< pwell >>
rect -2926 -2482 2926 2482
<< psubdiff >>
rect -2890 2412 -2794 2446
rect 2794 2412 2890 2446
rect -2890 2350 -2856 2412
rect 2856 2350 2890 2412
rect -2890 -2412 -2856 -2350
rect 2856 -2412 2890 -2350
rect -2890 -2446 -2794 -2412
rect 2794 -2446 2890 -2412
<< psubdiffcont >>
rect -2794 2412 2794 2446
rect -2890 -2350 -2856 2350
rect 2856 -2350 2890 2350
rect -2794 -2446 2794 -2412
<< xpolycontact >>
rect -2760 1884 -2622 2316
rect -2760 -2316 -2622 -1884
rect -2526 1884 -2388 2316
rect -2526 -2316 -2388 -1884
rect -2292 1884 -2154 2316
rect -2292 -2316 -2154 -1884
rect -2058 1884 -1920 2316
rect -2058 -2316 -1920 -1884
rect -1824 1884 -1686 2316
rect -1824 -2316 -1686 -1884
rect -1590 1884 -1452 2316
rect -1590 -2316 -1452 -1884
rect -1356 1884 -1218 2316
rect -1356 -2316 -1218 -1884
rect -1122 1884 -984 2316
rect -1122 -2316 -984 -1884
rect -888 1884 -750 2316
rect -888 -2316 -750 -1884
rect -654 1884 -516 2316
rect -654 -2316 -516 -1884
rect -420 1884 -282 2316
rect -420 -2316 -282 -1884
rect -186 1884 -48 2316
rect -186 -2316 -48 -1884
rect 48 1884 186 2316
rect 48 -2316 186 -1884
rect 282 1884 420 2316
rect 282 -2316 420 -1884
rect 516 1884 654 2316
rect 516 -2316 654 -1884
rect 750 1884 888 2316
rect 750 -2316 888 -1884
rect 984 1884 1122 2316
rect 984 -2316 1122 -1884
rect 1218 1884 1356 2316
rect 1218 -2316 1356 -1884
rect 1452 1884 1590 2316
rect 1452 -2316 1590 -1884
rect 1686 1884 1824 2316
rect 1686 -2316 1824 -1884
rect 1920 1884 2058 2316
rect 1920 -2316 2058 -1884
rect 2154 1884 2292 2316
rect 2154 -2316 2292 -1884
rect 2388 1884 2526 2316
rect 2388 -2316 2526 -1884
rect 2622 1884 2760 2316
rect 2622 -2316 2760 -1884
<< ppolyres >>
rect -2760 -1884 -2622 1884
rect -2526 -1884 -2388 1884
rect -2292 -1884 -2154 1884
rect -2058 -1884 -1920 1884
rect -1824 -1884 -1686 1884
rect -1590 -1884 -1452 1884
rect -1356 -1884 -1218 1884
rect -1122 -1884 -984 1884
rect -888 -1884 -750 1884
rect -654 -1884 -516 1884
rect -420 -1884 -282 1884
rect -186 -1884 -48 1884
rect 48 -1884 186 1884
rect 282 -1884 420 1884
rect 516 -1884 654 1884
rect 750 -1884 888 1884
rect 984 -1884 1122 1884
rect 1218 -1884 1356 1884
rect 1452 -1884 1590 1884
rect 1686 -1884 1824 1884
rect 1920 -1884 2058 1884
rect 2154 -1884 2292 1884
rect 2388 -1884 2526 1884
rect 2622 -1884 2760 1884
<< locali >>
rect -2890 2412 -2794 2446
rect 2794 2412 2890 2446
rect -2890 2350 -2856 2412
rect 2856 2350 2890 2412
rect -2890 -2412 -2856 -2350
rect 2856 -2412 2890 -2350
rect -2890 -2446 -2794 -2412
rect 2794 -2446 2890 -2412
<< viali >>
rect -2744 1901 -2638 2298
rect -2510 1901 -2404 2298
rect -2276 1901 -2170 2298
rect -2042 1901 -1936 2298
rect -1808 1901 -1702 2298
rect -1574 1901 -1468 2298
rect -1340 1901 -1234 2298
rect -1106 1901 -1000 2298
rect -872 1901 -766 2298
rect -638 1901 -532 2298
rect -404 1901 -298 2298
rect -170 1901 -64 2298
rect 64 1901 170 2298
rect 298 1901 404 2298
rect 532 1901 638 2298
rect 766 1901 872 2298
rect 1000 1901 1106 2298
rect 1234 1901 1340 2298
rect 1468 1901 1574 2298
rect 1702 1901 1808 2298
rect 1936 1901 2042 2298
rect 2170 1901 2276 2298
rect 2404 1901 2510 2298
rect 2638 1901 2744 2298
rect -2744 -2298 -2638 -1901
rect -2510 -2298 -2404 -1901
rect -2276 -2298 -2170 -1901
rect -2042 -2298 -1936 -1901
rect -1808 -2298 -1702 -1901
rect -1574 -2298 -1468 -1901
rect -1340 -2298 -1234 -1901
rect -1106 -2298 -1000 -1901
rect -872 -2298 -766 -1901
rect -638 -2298 -532 -1901
rect -404 -2298 -298 -1901
rect -170 -2298 -64 -1901
rect 64 -2298 170 -1901
rect 298 -2298 404 -1901
rect 532 -2298 638 -1901
rect 766 -2298 872 -1901
rect 1000 -2298 1106 -1901
rect 1234 -2298 1340 -1901
rect 1468 -2298 1574 -1901
rect 1702 -2298 1808 -1901
rect 1936 -2298 2042 -1901
rect 2170 -2298 2276 -1901
rect 2404 -2298 2510 -1901
rect 2638 -2298 2744 -1901
<< metal1 >>
rect -2750 2298 -2632 2310
rect -2750 1901 -2744 2298
rect -2638 1901 -2632 2298
rect -2750 1889 -2632 1901
rect -2516 2298 -2398 2310
rect -2516 1901 -2510 2298
rect -2404 1901 -2398 2298
rect -2516 1889 -2398 1901
rect -2282 2298 -2164 2310
rect -2282 1901 -2276 2298
rect -2170 1901 -2164 2298
rect -2282 1889 -2164 1901
rect -2048 2298 -1930 2310
rect -2048 1901 -2042 2298
rect -1936 1901 -1930 2298
rect -2048 1889 -1930 1901
rect -1814 2298 -1696 2310
rect -1814 1901 -1808 2298
rect -1702 1901 -1696 2298
rect -1814 1889 -1696 1901
rect -1580 2298 -1462 2310
rect -1580 1901 -1574 2298
rect -1468 1901 -1462 2298
rect -1580 1889 -1462 1901
rect -1346 2298 -1228 2310
rect -1346 1901 -1340 2298
rect -1234 1901 -1228 2298
rect -1346 1889 -1228 1901
rect -1112 2298 -994 2310
rect -1112 1901 -1106 2298
rect -1000 1901 -994 2298
rect -1112 1889 -994 1901
rect -878 2298 -760 2310
rect -878 1901 -872 2298
rect -766 1901 -760 2298
rect -878 1889 -760 1901
rect -644 2298 -526 2310
rect -644 1901 -638 2298
rect -532 1901 -526 2298
rect -644 1889 -526 1901
rect -410 2298 -292 2310
rect -410 1901 -404 2298
rect -298 1901 -292 2298
rect -410 1889 -292 1901
rect -176 2298 -58 2310
rect -176 1901 -170 2298
rect -64 1901 -58 2298
rect -176 1889 -58 1901
rect 58 2298 176 2310
rect 58 1901 64 2298
rect 170 1901 176 2298
rect 58 1889 176 1901
rect 292 2298 410 2310
rect 292 1901 298 2298
rect 404 1901 410 2298
rect 292 1889 410 1901
rect 526 2298 644 2310
rect 526 1901 532 2298
rect 638 1901 644 2298
rect 526 1889 644 1901
rect 760 2298 878 2310
rect 760 1901 766 2298
rect 872 1901 878 2298
rect 760 1889 878 1901
rect 994 2298 1112 2310
rect 994 1901 1000 2298
rect 1106 1901 1112 2298
rect 994 1889 1112 1901
rect 1228 2298 1346 2310
rect 1228 1901 1234 2298
rect 1340 1901 1346 2298
rect 1228 1889 1346 1901
rect 1462 2298 1580 2310
rect 1462 1901 1468 2298
rect 1574 1901 1580 2298
rect 1462 1889 1580 1901
rect 1696 2298 1814 2310
rect 1696 1901 1702 2298
rect 1808 1901 1814 2298
rect 1696 1889 1814 1901
rect 1930 2298 2048 2310
rect 1930 1901 1936 2298
rect 2042 1901 2048 2298
rect 1930 1889 2048 1901
rect 2164 2298 2282 2310
rect 2164 1901 2170 2298
rect 2276 1901 2282 2298
rect 2164 1889 2282 1901
rect 2398 2298 2516 2310
rect 2398 1901 2404 2298
rect 2510 1901 2516 2298
rect 2398 1889 2516 1901
rect 2632 2298 2750 2310
rect 2632 1901 2638 2298
rect 2744 1901 2750 2298
rect 2632 1889 2750 1901
rect -2750 -1901 -2632 -1889
rect -2750 -2298 -2744 -1901
rect -2638 -2298 -2632 -1901
rect -2750 -2310 -2632 -2298
rect -2516 -1901 -2398 -1889
rect -2516 -2298 -2510 -1901
rect -2404 -2298 -2398 -1901
rect -2516 -2310 -2398 -2298
rect -2282 -1901 -2164 -1889
rect -2282 -2298 -2276 -1901
rect -2170 -2298 -2164 -1901
rect -2282 -2310 -2164 -2298
rect -2048 -1901 -1930 -1889
rect -2048 -2298 -2042 -1901
rect -1936 -2298 -1930 -1901
rect -2048 -2310 -1930 -2298
rect -1814 -1901 -1696 -1889
rect -1814 -2298 -1808 -1901
rect -1702 -2298 -1696 -1901
rect -1814 -2310 -1696 -2298
rect -1580 -1901 -1462 -1889
rect -1580 -2298 -1574 -1901
rect -1468 -2298 -1462 -1901
rect -1580 -2310 -1462 -2298
rect -1346 -1901 -1228 -1889
rect -1346 -2298 -1340 -1901
rect -1234 -2298 -1228 -1901
rect -1346 -2310 -1228 -2298
rect -1112 -1901 -994 -1889
rect -1112 -2298 -1106 -1901
rect -1000 -2298 -994 -1901
rect -1112 -2310 -994 -2298
rect -878 -1901 -760 -1889
rect -878 -2298 -872 -1901
rect -766 -2298 -760 -1901
rect -878 -2310 -760 -2298
rect -644 -1901 -526 -1889
rect -644 -2298 -638 -1901
rect -532 -2298 -526 -1901
rect -644 -2310 -526 -2298
rect -410 -1901 -292 -1889
rect -410 -2298 -404 -1901
rect -298 -2298 -292 -1901
rect -410 -2310 -292 -2298
rect -176 -1901 -58 -1889
rect -176 -2298 -170 -1901
rect -64 -2298 -58 -1901
rect -176 -2310 -58 -2298
rect 58 -1901 176 -1889
rect 58 -2298 64 -1901
rect 170 -2298 176 -1901
rect 58 -2310 176 -2298
rect 292 -1901 410 -1889
rect 292 -2298 298 -1901
rect 404 -2298 410 -1901
rect 292 -2310 410 -2298
rect 526 -1901 644 -1889
rect 526 -2298 532 -1901
rect 638 -2298 644 -1901
rect 526 -2310 644 -2298
rect 760 -1901 878 -1889
rect 760 -2298 766 -1901
rect 872 -2298 878 -1901
rect 760 -2310 878 -2298
rect 994 -1901 1112 -1889
rect 994 -2298 1000 -1901
rect 1106 -2298 1112 -1901
rect 994 -2310 1112 -2298
rect 1228 -1901 1346 -1889
rect 1228 -2298 1234 -1901
rect 1340 -2298 1346 -1901
rect 1228 -2310 1346 -2298
rect 1462 -1901 1580 -1889
rect 1462 -2298 1468 -1901
rect 1574 -2298 1580 -1901
rect 1462 -2310 1580 -2298
rect 1696 -1901 1814 -1889
rect 1696 -2298 1702 -1901
rect 1808 -2298 1814 -1901
rect 1696 -2310 1814 -2298
rect 1930 -1901 2048 -1889
rect 1930 -2298 1936 -1901
rect 2042 -2298 2048 -1901
rect 1930 -2310 2048 -2298
rect 2164 -1901 2282 -1889
rect 2164 -2298 2170 -1901
rect 2276 -2298 2282 -1901
rect 2164 -2310 2282 -2298
rect 2398 -1901 2516 -1889
rect 2398 -2298 2404 -1901
rect 2510 -2298 2516 -1901
rect 2398 -2310 2516 -2298
rect 2632 -1901 2750 -1889
rect 2632 -2298 2638 -1901
rect 2744 -2298 2750 -1901
rect 2632 -2310 2750 -2298
<< properties >>
string FIXED_BBOX -2873 -2429 2873 2429
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.690 l 19.0 m 1 nx 24 wmin 0.690 lmin 0.50 rho 319.8 val 9.37k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
