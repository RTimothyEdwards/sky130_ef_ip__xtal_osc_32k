VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_ip__xtal_osc_32k
  CLASS BLOCK ;
  FOREIGN sky130_ef_ip__xtal_osc_32k ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.170 BY 132.790 ;
  PIN in
    ANTENNAGATEAREA 0.420000 ;
    ANTENNADIFFAREA 0.526800 ;
    PORT
      LAYER met1 ;
        RECT 0.000 130.895 1.000 131.895 ;
    END
  END in
  PIN out
    PORT
      LAYER met1 ;
        RECT 0.000 55.045 1.000 56.045 ;
    END
  END out
  PIN avdd
    ANTENNADIFFAREA 200.228592 ;
    PORT
      LAYER met2 ;
        RECT 0.000 84.540 1.710 104.540 ;
    END
    PORT
      LAYER met2 ;
        RECT 68.460 84.540 70.170 104.540 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.000 7.240 1.710 27.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 68.460 7.240 70.170 27.240 ;
    END
  END avdd
  PIN avss
    ANTENNADIFFAREA 172.646790 ;
    PORT
      LAYER met2 ;
        RECT 0.000 28.780 1.840 48.780 ;
    END
    PORT
      LAYER met2 ;
        RECT 68.330 28.780 70.170 48.780 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.000 105.965 2.075 125.965 ;
    END
    PORT
      LAYER met2 ;
        RECT 68.240 105.965 70.170 125.965 ;
    END
  END avss
  PIN dvss
    ANTENNADIFFAREA 15.428800 ;
    PORT
      LAYER met2 ;
        RECT 67.735 74.670 70.170 75.670 ;
    END
  END dvss
  PIN dvdd
    ANTENNADIFFAREA 4.959600 ;
    PORT
      LAYER met2 ;
        RECT 67.885 62.295 70.170 63.295 ;
    END
  END dvdd
  PIN ena
    ANTENNAGATEAREA 0.585000 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met2 ;
        RECT 69.170 72.285 70.170 73.285 ;
    END
  END ena
  PIN dout
    PORT
      LAYER met1 ;
        RECT 69.170 76.485 70.170 77.485 ;
    END
  END dout
  PIN boost
    ANTENNAGATEAREA 0.510000 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met2 ;
        RECT 69.170 59.870 70.170 60.870 ;
    END
  END boost
  OBS
      LAYER nwell ;
        RECT 0.000 131.210 70.170 132.790 ;
        RECT 0.000 1.730 1.580 131.210 ;
        RECT 0.000 0.000 70.170 1.730 ;
      LAYER li1 ;
        RECT 0.285 0.340 70.040 132.460 ;
      LAYER met1 ;
        RECT 0.070 132.175 70.135 132.720 ;
        RECT 1.280 130.615 70.135 132.175 ;
        RECT 0.070 77.765 70.135 130.615 ;
        RECT 0.070 76.205 68.890 77.765 ;
        RECT 0.070 56.325 70.135 76.205 ;
        RECT 1.280 54.765 70.135 56.325 ;
        RECT 0.070 0.080 70.135 54.765 ;
      LAYER met2 ;
        RECT 2.355 105.685 67.960 125.970 ;
        RECT 0.335 104.820 69.170 105.685 ;
        RECT 1.990 84.260 68.180 104.820 ;
        RECT 0.335 75.950 69.170 84.260 ;
        RECT 0.335 74.390 67.455 75.950 ;
        RECT 0.335 73.565 69.170 74.390 ;
        RECT 0.335 72.005 68.890 73.565 ;
        RECT 0.335 63.575 69.170 72.005 ;
        RECT 0.335 62.015 67.605 63.575 ;
        RECT 0.335 61.150 69.170 62.015 ;
        RECT 0.335 59.590 68.890 61.150 ;
        RECT 0.335 49.060 69.170 59.590 ;
        RECT 2.120 28.500 68.050 49.060 ;
        RECT 0.335 27.520 69.170 28.500 ;
        RECT 1.990 7.240 68.180 27.520 ;
  END
END sky130_ef_ip__xtal_osc_32k
END LIBRARY

