magic
tech sky130A
magscale 1 2
timestamp 1699546087
<< dnwell >>
rect 110 15744 13924 26448
rect 110 10806 12214 15744
rect 110 110 13924 10806
<< nwell >>
rect 0 26242 14034 26558
rect 0 346 316 26242
rect 13718 15952 14034 26242
rect 12008 15636 14034 15952
rect 6834 14118 7450 14726
rect 9914 14118 10006 14726
rect 12008 14704 12324 15636
rect 6834 14048 10006 14118
rect 9914 13440 10006 14048
rect 11980 13358 12324 14704
rect 13536 13858 13622 14426
rect 10754 13134 12324 13358
rect 11980 11797 12324 13134
rect 12008 10916 12324 11797
rect 12008 10600 14034 10916
rect 13718 346 14034 10600
rect 0 0 14034 346
<< mvnsubdiff >>
rect 67 26471 13967 26491
rect 67 26437 147 26471
rect 13887 26437 13967 26471
rect 67 26417 13967 26437
rect 67 26411 141 26417
rect 67 147 87 26411
rect 121 147 141 26411
rect 13893 26411 13967 26417
rect 13893 15798 13913 26411
rect 13947 15798 13967 26411
rect 13893 15779 13967 15798
rect 12173 15759 13967 15779
rect 12173 15725 12267 15759
rect 13897 15725 13967 15759
rect 12173 15709 13967 15725
rect 12173 10833 12193 15709
rect 12227 15705 13967 15709
rect 12227 10837 12247 15705
rect 12227 10833 13967 10837
rect 12173 10817 13967 10833
rect 12173 10783 12263 10817
rect 13877 10783 13967 10817
rect 12173 10763 13967 10783
rect 67 141 141 147
rect 13893 10748 13967 10763
rect 13893 150 13913 10748
rect 13947 150 13967 10748
rect 13893 141 13967 150
rect 67 121 13967 141
rect 67 87 147 121
rect 13887 87 13967 121
rect 67 67 13967 87
<< mvnsubdiffcont >>
rect 147 26437 13887 26471
rect 87 147 121 26411
rect 13913 15798 13947 26411
rect 12267 15725 13897 15759
rect 12193 10833 12227 15709
rect 12263 10783 13877 10817
rect 13913 150 13947 10748
rect 147 87 13887 121
<< locali >>
rect 87 26437 147 26471
rect 13887 26437 13947 26471
rect 87 26411 121 26437
rect 13913 26411 13947 26437
rect 9295 16053 9546 16055
rect 9014 16034 9546 16053
rect 9014 15751 10050 16034
rect 13913 15759 13947 15798
rect 9014 15610 9546 15751
rect 12193 15725 12267 15759
rect 13897 15725 13947 15759
rect 12193 15709 12227 15725
rect 9286 15359 9546 15610
rect 9304 15261 9546 15359
rect 9286 15260 9546 15261
rect 9397 15224 9546 15260
rect 9397 15156 9531 15224
rect 6919 14648 9936 14809
rect 6919 14226 7534 14648
rect 7973 14226 8153 14648
rect 8592 14226 8772 14648
rect 9201 14226 9381 14648
rect 9810 14226 9936 14648
rect 6919 14200 9936 14226
rect 6919 14199 8254 14200
rect 6919 14198 7613 14199
rect 6919 14117 6975 14198
rect 7481 14117 7613 14198
rect 6919 13972 7613 14117
rect 7688 13973 8254 14199
rect 8329 14199 9936 14200
rect 8329 13973 8855 14199
rect 7688 13972 8855 13973
rect 8930 14197 9936 14199
rect 8930 13972 9683 14197
rect 6919 13970 9683 13972
rect 9758 13970 9936 14197
rect 6919 13950 9936 13970
rect 7350 13540 7539 13950
rect 7973 13540 8162 13950
rect 8578 13540 8767 13950
rect 9206 13540 9395 13950
rect 9810 13540 9936 13950
rect 6908 13419 9936 13540
rect 6811 13155 10052 13274
rect 7249 12761 7385 13155
rect 7811 12761 7955 13155
rect 8359 12761 8503 13155
rect 8929 12761 9073 13155
rect 9482 12761 9626 13155
rect 6810 12741 10051 12761
rect 6810 12738 8751 12741
rect 6810 12737 7645 12738
rect 6810 12567 7074 12737
rect 7240 12568 7645 12737
rect 7811 12568 8195 12738
rect 8361 12571 8751 12738
rect 8917 12571 9309 12741
rect 9475 12738 10051 12741
rect 9475 12571 9808 12738
rect 8361 12568 9808 12571
rect 9974 12568 10051 12738
rect 7240 12567 10051 12568
rect 6810 12563 10051 12567
rect 7254 12160 7394 12563
rect 7806 12160 7950 12563
rect 8363 12160 8507 12563
rect 8921 12160 9065 12563
rect 9478 12160 9622 12563
rect 6805 12077 10054 12160
rect 6805 12073 8541 12077
rect 6805 12003 8147 12073
rect 6805 11899 6894 12003
rect 7913 11903 8147 12003
rect 8313 11907 8541 12073
rect 8707 12065 10054 12077
rect 8707 11907 9294 12065
rect 8313 11903 9294 11907
rect 7913 11899 9294 11903
rect 6805 11895 9294 11899
rect 9460 11895 10054 12065
rect 6805 11823 10054 11895
rect 8361 11406 8506 11823
rect 8916 11409 9060 11823
rect 9482 11409 9626 11823
rect 13484 14919 13931 15021
rect 13494 14898 13931 14919
rect 12860 14704 12992 14784
rect 12860 11798 12907 14704
rect 12966 11798 12992 14704
rect 13494 14638 13650 14898
rect 13492 13894 13671 14390
rect 13573 13199 13661 13583
rect 13235 13197 14008 13199
rect 13234 13190 14008 13197
rect 13234 13132 13252 13190
rect 13805 13132 14008 13190
rect 13234 13127 14008 13132
rect 13235 13124 14008 13127
rect 12860 11694 12992 11798
rect 12668 11444 13024 11456
rect 12668 11264 12850 11444
rect 13012 11264 13024 11444
rect 12668 11253 13024 11264
rect 12193 10817 12227 10833
rect 12193 10783 12263 10817
rect 13877 10783 13947 10817
rect 13913 10748 13947 10783
rect 87 121 121 147
rect 13913 121 13947 150
rect 87 87 147 121
rect 13887 87 13947 121
<< viali >>
rect 631 26471 13767 26492
rect 631 26437 13767 26471
rect 631 26426 13767 26437
rect 13892 25551 13913 25982
rect 13913 25551 13947 25982
rect 13947 25551 13967 25982
rect 57 21094 87 25178
rect 87 21094 121 25178
rect 121 21094 141 25178
rect 423 21221 458 25184
rect 10008 21202 10060 25165
rect 10311 21202 10363 25165
rect 13596 21207 13648 25170
rect 13895 21204 13913 25186
rect 13913 21204 13947 25186
rect 13947 21204 13969 25186
rect 66 16924 87 20888
rect 87 16924 121 20888
rect 121 16924 141 20888
rect 13893 16918 13913 20884
rect 13913 16918 13947 20884
rect 13947 16918 13967 20884
rect 57 11451 87 16777
rect 87 11451 121 16777
rect 121 11451 144 16777
rect 13891 15837 13913 16768
rect 13913 15837 13947 16768
rect 13947 15837 13966 16768
rect 12373 15759 13839 15776
rect 12373 15725 13839 15759
rect 12373 15712 13839 15725
rect 507 11356 580 15488
rect 9014 15261 9304 15359
rect 9668 15278 9962 15360
rect 9531 15156 10099 15224
rect 6975 14117 7481 14198
rect 7613 13972 7688 14199
rect 8254 13973 8329 14200
rect 8855 13972 8930 14199
rect 9683 13970 9758 14197
rect 7074 12567 7240 12737
rect 7645 12568 7811 12738
rect 8195 12568 8361 12738
rect 8751 12571 8917 12741
rect 9309 12571 9475 12741
rect 9808 12568 9974 12738
rect 6894 11899 7913 12003
rect 8147 11903 8313 12073
rect 8541 11907 8707 12077
rect 9294 11895 9460 12065
rect 12180 10864 12193 15671
rect 12193 10864 12227 15671
rect 12227 10864 12240 15671
rect 12907 11798 12966 14704
rect 13252 13132 13805 13190
rect 12850 11264 13012 11444
rect 12341 10817 13778 10836
rect 12341 10783 13778 10817
rect 12341 10778 13778 10783
rect 368 5766 420 9742
rect 13614 5764 13666 9740
rect 13887 5776 13913 10643
rect 13913 5776 13947 10643
rect 13947 5776 13950 10643
rect 67 1459 87 5440
rect 87 1459 121 5440
rect 121 1459 142 5440
rect 13894 1462 13913 5428
rect 13913 1462 13947 5428
rect 13947 1462 13967 5428
rect 66 584 87 1014
rect 87 584 121 1014
rect 121 584 141 1014
rect 175 121 13853 144
rect 175 87 13853 121
rect 175 68 13853 87
<< metal1 >>
rect 13806 26543 14027 26544
rect 512 26492 14027 26543
rect 512 26426 631 26492
rect 13767 26426 14027 26492
rect 512 26396 14027 26426
rect 0 26328 200 26379
rect 0 26241 10224 26328
rect 0 26179 200 26241
rect 10137 25992 10224 26241
rect 554 25560 790 25992
rect 886 25560 1122 25992
rect 1218 25560 1454 25992
rect 1550 25560 1786 25992
rect 1882 25560 2118 25992
rect 2214 25560 2450 25992
rect 2546 25560 2782 25992
rect 2878 25560 3114 25992
rect 3210 25560 3446 25992
rect 3542 25560 3778 25992
rect 3874 25560 4110 25992
rect 4206 25560 4442 25992
rect 4538 25560 4774 25992
rect 4870 25560 5106 25992
rect 5202 25560 5438 25992
rect 5534 25560 5770 25992
rect 5866 25560 6102 25992
rect 6198 25560 6434 25992
rect 6530 25560 6766 25992
rect 6862 25560 7098 25992
rect 7194 25560 7430 25992
rect 7526 25560 7762 25992
rect 7858 25560 8094 25992
rect 8190 25560 8426 25992
rect 8522 25560 8758 25992
rect 8854 25560 9090 25992
rect 9186 25560 9422 25992
rect 9518 25560 9754 25992
rect 9850 25560 10224 25992
rect 13806 25982 14027 26396
rect 14 25178 178 25213
rect 417 25184 464 25196
rect 14 21094 57 25178
rect 141 21094 178 25178
rect 405 21221 415 25184
rect 467 21221 477 25184
rect 10002 25165 10066 25177
rect 417 21209 464 21221
rect 9998 21202 10008 25165
rect 10060 21202 10070 25165
rect 10002 21190 10066 21202
rect 14 20888 178 21094
rect 14 16924 66 20888
rect 141 16924 178 20888
rect 14 16777 178 16924
rect 14 11451 57 16777
rect 144 11451 178 16777
rect 554 15925 624 16592
rect 720 16160 956 16592
rect 1052 16160 1288 16592
rect 1384 16160 1620 16592
rect 1716 16160 1952 16592
rect 2048 16160 2284 16592
rect 2380 16160 2616 16592
rect 2712 16160 2948 16592
rect 3044 16160 3280 16592
rect 3376 16160 3612 16592
rect 3708 16160 3944 16592
rect 4040 16160 4276 16592
rect 4372 16160 4608 16592
rect 4704 16160 4940 16592
rect 5036 16160 5272 16592
rect 5368 16160 5604 16592
rect 5700 16160 5936 16592
rect 6032 16160 6268 16592
rect 6364 16160 6600 16592
rect 6696 16160 6932 16592
rect 7028 16160 7264 16592
rect 7360 16160 7596 16592
rect 7692 16160 7928 16592
rect 8024 16160 8260 16592
rect 8356 16160 8592 16592
rect 8688 16160 8924 16592
rect 9020 16160 9256 16592
rect 9352 16160 9588 16592
rect 9684 16160 9920 16592
rect 554 15826 6484 15925
rect 501 15488 586 15500
rect 14 11411 178 11451
rect 497 11356 507 15488
rect 580 11356 590 15488
rect 670 15148 1042 15580
rect 1138 15148 1510 15580
rect 1606 15148 1978 15580
rect 2074 15148 2446 15580
rect 2542 15148 2914 15580
rect 3010 15148 3382 15580
rect 3478 15148 3850 15580
rect 3946 15148 4318 15580
rect 4414 15148 4786 15580
rect 4882 15148 5254 15580
rect 5350 15148 5722 15580
rect 5818 15148 6190 15580
rect 6387 14071 6484 15826
rect 10137 15506 10224 25560
rect 10450 25550 10686 25982
rect 10782 25550 11018 25982
rect 11114 25550 11350 25982
rect 11446 25550 11682 25982
rect 11778 25550 12014 25982
rect 12110 25550 12346 25982
rect 12442 25550 12678 25982
rect 12774 25550 13010 25982
rect 13106 25550 13342 25982
rect 13438 25551 13892 25982
rect 13967 25551 14027 25982
rect 13438 25550 14027 25551
rect 13806 25186 14027 25550
rect 10305 25165 10369 25177
rect 13590 25170 13654 25182
rect 10301 21202 10311 25165
rect 10363 21202 10373 25165
rect 13586 21207 13596 25170
rect 13648 21207 13658 25170
rect 10305 21190 10369 21202
rect 13590 21195 13654 21207
rect 13806 21204 13895 25186
rect 13969 21204 14027 25186
rect 13806 20884 14027 21204
rect 13806 16918 13893 20884
rect 13967 16918 14027 20884
rect 13806 16768 14027 16918
rect 9107 15438 10224 15506
rect 10332 16171 10504 16236
rect 9107 15437 10214 15438
rect 9002 15359 9316 15365
rect 9002 15261 9014 15359
rect 9304 15261 9316 15359
rect 9656 15360 9974 15366
rect 9656 15278 9668 15360
rect 9962 15278 9974 15360
rect 9656 15272 9974 15278
rect 9002 15255 9316 15261
rect 9023 15046 9284 15255
rect 9519 15224 10111 15230
rect 9519 15156 9531 15224
rect 10099 15156 10111 15224
rect 9519 15150 10111 15156
rect 9610 15046 9984 15150
rect 9023 14829 9977 15046
rect 9023 14828 9284 14829
rect 9967 14828 9977 14829
rect 10045 14828 10055 15046
rect 10003 14644 10071 14654
rect 8992 14532 9416 14533
rect 7706 14481 9416 14532
rect 9562 14486 10003 14528
rect 7706 14480 9042 14481
rect 7629 14215 7675 14428
rect 6963 14198 7493 14204
rect 6963 14117 6975 14198
rect 7481 14117 7493 14198
rect 6963 14111 7493 14117
rect 7466 14071 7510 14073
rect 6387 14027 7510 14071
rect 6387 12163 6484 14027
rect 6921 13758 7076 13802
rect 6921 13616 6965 13758
rect 7030 13651 7193 13692
rect 6892 13432 6902 13616
rect 6967 13432 6977 13616
rect 6911 13426 6965 13432
rect 6646 13168 6656 13326
rect 6715 13168 6725 13326
rect 6662 12286 6711 13168
rect 6911 12876 6954 13426
rect 7030 13418 7071 13651
rect 7021 13260 7031 13418
rect 7090 13260 7100 13418
rect 7229 13264 7304 13825
rect 7466 13803 7510 14027
rect 7571 13979 7581 14215
rect 7744 13979 7754 14215
rect 7607 13972 7613 13979
rect 7688 13972 7694 13979
rect 7607 13960 7694 13972
rect 7466 13759 7686 13803
rect 7030 13254 7071 13260
rect 7183 13103 7193 13264
rect 7350 13103 7360 13264
rect 6999 13023 7340 13045
rect 6999 13004 7291 13023
rect 7129 12846 7179 12965
rect 7281 12856 7291 13004
rect 7348 12856 7358 13023
rect 7466 12884 7510 13759
rect 7850 13736 7891 14424
rect 8270 14212 8316 14427
rect 8248 14210 8335 14212
rect 8202 13974 8212 14210
rect 8375 13974 8385 14210
rect 8248 13973 8254 13974
rect 8329 13973 8335 13974
rect 8248 13961 8335 13973
rect 7734 13516 7775 13683
rect 8247 13516 8291 13826
rect 8476 13736 8517 14424
rect 8867 14211 8913 14425
rect 8849 14202 8936 14211
rect 8805 13966 8815 14202
rect 8978 13966 8988 14202
rect 8849 13960 8936 13966
rect 7734 13472 8291 13516
rect 8358 13511 8399 13685
rect 8847 13511 8891 13825
rect 9075 13739 9116 14427
rect 9364 14408 9416 14481
rect 10003 14457 10071 14467
rect 9364 14360 9547 14408
rect 9364 13801 9416 14360
rect 9699 14209 9748 14424
rect 10143 14371 10197 15437
rect 10332 15354 10397 16171
rect 10616 16150 10852 16582
rect 10948 16150 11184 16582
rect 11280 16150 11516 16582
rect 11612 16150 11848 16582
rect 11944 16150 12180 16582
rect 12276 16150 12512 16582
rect 12608 16150 12844 16582
rect 12940 16150 13176 16582
rect 13272 16150 13508 16582
rect 13806 15892 13891 16768
rect 12116 15837 13891 15892
rect 13966 15837 14027 16768
rect 12116 15776 14027 15837
rect 12116 15712 12373 15776
rect 13839 15712 14027 15776
rect 12116 15671 14027 15712
rect 10536 15492 10546 15650
rect 11992 15492 12002 15650
rect 9951 14317 10197 14371
rect 10272 15238 10397 15354
rect 9677 14204 9764 14209
rect 9629 13968 9639 14204
rect 9802 13968 9812 14204
rect 9677 13958 9764 13968
rect 9364 13757 9540 13801
rect 9364 13752 9528 13757
rect 7734 13424 7775 13472
rect 7579 13366 7589 13424
rect 7775 13366 7785 13424
rect 7587 13012 7628 13366
rect 7684 12846 7734 12966
rect 8037 12886 8081 13472
rect 8358 13467 8891 13511
rect 8358 13416 8399 13467
rect 8139 13375 8399 13416
rect 8139 13015 8180 13375
rect 6909 12796 7179 12846
rect 7459 12796 7734 12846
rect 8233 12843 8283 12967
rect 8591 12876 8635 13467
rect 8970 13392 9011 13683
rect 9364 13679 9416 13752
rect 9699 13731 9748 13958
rect 9364 13627 9657 13679
rect 8970 13381 9047 13392
rect 8702 13340 9047 13381
rect 8702 13015 8743 13340
rect 8973 13329 9047 13340
rect 9270 13329 9280 13392
rect 8792 12843 8842 12963
rect 6909 12339 6959 12796
rect 7068 12737 7246 12749
rect 7068 12567 7074 12737
rect 7240 12567 7246 12737
rect 7068 12555 7246 12567
rect 7131 12344 7183 12555
rect 7459 12339 7509 12796
rect 8019 12793 8283 12843
rect 8583 12793 8842 12843
rect 7639 12738 7817 12750
rect 7639 12568 7645 12738
rect 7811 12568 7817 12738
rect 7639 12556 7817 12568
rect 7695 12342 7747 12556
rect 8019 12340 8069 12793
rect 8189 12738 8367 12750
rect 8189 12568 8195 12738
rect 8361 12568 8367 12738
rect 8189 12556 8367 12568
rect 8249 12340 8301 12556
rect 8583 12340 8633 12793
rect 8745 12741 8923 12753
rect 8745 12571 8751 12741
rect 8917 12571 8923 12741
rect 8745 12559 8923 12571
rect 8803 12338 8855 12559
rect 8973 12535 9014 13329
rect 9364 13206 9416 13627
rect 9505 13327 9515 13390
rect 9738 13385 9748 13390
rect 9951 13385 10005 14317
rect 10272 14086 10337 15238
rect 10379 14438 10389 14615
rect 10457 14498 10467 14615
rect 10768 14554 11210 14615
rect 10768 14498 10829 14554
rect 10457 14438 10829 14498
rect 10396 14437 10829 14438
rect 10202 14015 10337 14086
rect 10399 14098 10548 14160
rect 10054 13596 10064 13868
rect 10139 13596 10149 13868
rect 9738 13331 10005 13385
rect 9738 13327 9748 13331
rect 9123 13154 9416 13206
rect 9123 12888 9175 13154
rect 10073 13061 10127 13596
rect 9224 13031 10127 13061
rect 9224 13007 9522 13031
rect 9339 12843 9389 12959
rect 9512 12864 9522 13007
rect 9579 13007 10127 13031
rect 9579 12864 9589 13007
rect 9127 12793 9389 12843
rect 8952 12358 8962 12535
rect 9033 12358 9043 12535
rect 9127 12338 9177 12793
rect 9303 12741 9481 12753
rect 9303 12571 9309 12741
rect 9475 12571 9481 12741
rect 9303 12559 9481 12571
rect 9364 12347 9416 12559
rect 6662 12237 7086 12286
rect 9684 12283 9741 12965
rect 10202 12955 10267 14015
rect 9889 12893 10127 12953
rect 9802 12738 9980 12750
rect 9802 12568 9808 12738
rect 9974 12568 9980 12738
rect 9802 12556 9980 12568
rect 9913 12340 9973 12556
rect 7554 12225 9857 12283
rect 6387 12124 8072 12163
rect 501 11344 586 11356
rect 0 11166 200 11209
rect 0 11059 686 11166
rect 0 11009 200 11059
rect 904 10948 1276 11380
rect 1372 10948 1744 11380
rect 1840 10948 2212 11380
rect 2308 10948 2680 11380
rect 2776 10948 3148 11380
rect 3244 10948 3616 11380
rect 3712 10948 4084 11380
rect 4180 10948 4552 11380
rect 4648 10948 5020 11380
rect 5116 10948 5488 11380
rect 5584 10948 5956 11380
rect 6387 11214 6484 12124
rect 6882 12003 7925 12009
rect 6882 11899 6894 12003
rect 7913 11899 7925 12003
rect 6882 11893 7925 11899
rect 8033 11613 8072 12124
rect 8141 12073 8319 12085
rect 8535 12077 8713 12089
rect 8137 11903 8147 12073
rect 8313 11903 8323 12073
rect 8531 11907 8541 12077
rect 8707 11907 8717 12077
rect 8953 11907 8963 12084
rect 9034 11907 9044 12084
rect 8141 11891 8319 11903
rect 8535 11895 8713 11907
rect 8248 11611 8300 11891
rect 8581 11613 8633 11895
rect 8964 11688 9012 11907
rect 8792 11640 9012 11688
rect 9144 11621 9188 12225
rect 9288 12065 9466 12077
rect 9284 11895 9294 12065
rect 9460 11895 9470 12065
rect 9288 11883 9466 11895
rect 9346 11615 9398 11883
rect 9702 11625 9757 12225
rect 9792 11929 9800 11997
rect 10000 11929 10010 11997
rect 9909 11620 9959 11929
rect 8106 11561 9672 11568
rect 8106 11512 9607 11561
rect 9597 11384 9607 11512
rect 9678 11384 9688 11561
rect 9616 11377 9672 11384
rect 9802 11337 9854 11570
rect 9792 11269 9802 11337
rect 10002 11269 10012 11337
rect 6171 11092 6484 11214
rect 10067 10672 10127 12893
rect 10182 12901 10267 12955
rect 10182 12004 10247 12901
rect 10399 12849 10461 14098
rect 10507 13659 10701 13664
rect 10503 13461 10513 13659
rect 10695 13461 10705 13659
rect 12116 13586 12180 15671
rect 10295 12789 10461 12849
rect 10507 13036 10701 13461
rect 10507 12844 10518 13036
rect 10697 12844 10707 13036
rect 11968 12910 12180 13586
rect 10507 12835 10701 12844
rect 10167 11992 10258 12004
rect 10167 11815 10177 11992
rect 10248 11815 10258 11992
rect 10295 11721 10355 12789
rect 10195 11661 10355 11721
rect 10404 12578 10559 12638
rect 10195 11605 10255 11661
rect 10177 11428 10187 11605
rect 10258 11428 10268 11605
rect 10404 11334 10464 12578
rect 10222 11266 10232 11334
rect 10432 11267 10464 11334
rect 10432 11266 10442 11267
rect 10544 10833 10554 10994
rect 11980 10833 11990 10994
rect 12116 10864 12180 12910
rect 12240 10911 12341 15671
rect 13834 15442 14034 15497
rect 12647 15365 14034 15442
rect 12647 14542 12724 15365
rect 13834 15297 14034 15365
rect 12838 15118 13568 15136
rect 12838 14948 13382 15118
rect 13547 14948 13568 15118
rect 12838 14934 13568 14948
rect 12838 14704 13058 14934
rect 12451 11864 12461 11918
rect 12576 11864 12586 11918
rect 12524 11290 12576 11864
rect 12636 11150 12734 11852
rect 12838 11798 12907 14704
rect 12966 13407 13058 14704
rect 13596 14752 13820 14801
rect 13596 14523 13645 14752
rect 13580 14466 13590 14523
rect 13649 14466 13660 14523
rect 13712 13930 13765 14274
rect 13594 13730 13765 13930
rect 13805 13669 13845 14003
rect 13388 13629 13845 13669
rect 13088 13438 13098 13490
rect 13188 13489 13198 13490
rect 13388 13489 13430 13629
rect 13188 13479 13430 13489
rect 13188 13449 13392 13479
rect 13188 13438 13198 13449
rect 13590 13447 13600 13499
rect 13652 13487 13662 13499
rect 13652 13447 13849 13487
rect 12966 13315 13377 13407
rect 13464 13346 13789 13391
rect 12966 13198 13146 13315
rect 12966 13190 13818 13198
rect 12966 13132 13252 13190
rect 13805 13132 13818 13190
rect 12966 13122 13818 13132
rect 12966 12951 13146 13122
rect 13465 12979 13475 13034
rect 13529 13024 13539 13034
rect 13529 12990 13847 13024
rect 13529 12979 13539 12990
rect 12966 12864 13800 12951
rect 12966 11798 13058 12864
rect 13882 12828 13981 14281
rect 13667 12730 13981 12828
rect 12838 11485 13058 11798
rect 12838 11444 13566 11485
rect 12838 11264 12850 11444
rect 13012 11264 13566 11444
rect 12838 11253 13566 11264
rect 13667 11150 13765 12730
rect 12636 11052 13765 11150
rect 12240 10864 14004 10911
rect 12116 10836 14004 10864
rect 12116 10778 12341 10836
rect 13778 10778 14004 10836
rect 12116 10770 14004 10778
rect 12117 10760 14004 10770
rect 10067 10612 13528 10672
rect 510 9982 747 10414
rect 841 9982 1078 10414
rect 1172 9982 1409 10414
rect 1503 9982 1740 10414
rect 1834 9982 2071 10414
rect 2165 9982 2402 10414
rect 2496 9982 2733 10414
rect 2827 9982 3064 10414
rect 3158 9982 3395 10414
rect 3489 9982 3726 10414
rect 3820 9982 4057 10414
rect 4151 9982 4388 10414
rect 4482 9982 4719 10414
rect 4813 9982 5050 10414
rect 5144 9982 5381 10414
rect 5475 9982 5712 10414
rect 5806 9982 6043 10414
rect 6137 9982 6374 10414
rect 6468 9982 6705 10414
rect 6799 9982 7036 10414
rect 7130 9982 7367 10414
rect 7461 9982 7698 10414
rect 7792 9982 8029 10414
rect 8123 9982 8360 10414
rect 8454 9982 8691 10414
rect 8785 9982 9022 10414
rect 9116 9982 9353 10414
rect 9447 9982 9684 10414
rect 9778 9982 10015 10414
rect 10109 9982 10346 10414
rect 10440 9982 10677 10414
rect 10771 9982 11008 10414
rect 11102 9982 11339 10414
rect 11433 9982 11670 10414
rect 11764 9982 12001 10414
rect 12095 9982 12332 10414
rect 12426 9982 12663 10414
rect 12757 9982 12994 10414
rect 13088 9982 13325 10414
rect 13458 9982 13528 10612
rect 13853 10643 14004 10760
rect 362 9742 426 9754
rect 358 5766 368 9742
rect 420 5766 430 9742
rect 13608 9740 13672 9752
rect 362 5754 426 5766
rect 13604 5764 13614 9740
rect 13666 5764 13676 9740
rect 13853 5776 13887 10643
rect 13950 5776 14004 10643
rect 13608 5752 13672 5764
rect 61 5440 148 5452
rect 57 1459 67 5440
rect 142 1459 152 5440
rect 13853 5428 14004 5776
rect 13853 1462 13894 5428
rect 13967 1462 14004 5428
rect 60 1447 148 1459
rect 60 1014 147 1447
rect 60 584 66 1014
rect 141 584 580 1014
rect 60 582 580 584
rect 676 582 912 1014
rect 1008 582 1244 1014
rect 1340 582 1576 1014
rect 1672 582 1908 1014
rect 2004 582 2240 1014
rect 2336 582 2572 1014
rect 2668 582 2904 1014
rect 3000 582 3236 1014
rect 3332 582 3568 1014
rect 3664 582 3900 1014
rect 3996 582 4232 1014
rect 4328 582 4564 1014
rect 4660 582 4896 1014
rect 4992 582 5228 1014
rect 5324 582 5560 1014
rect 5656 582 5892 1014
rect 5988 582 6224 1014
rect 6320 582 6556 1014
rect 6652 582 6888 1014
rect 6984 582 7220 1014
rect 7316 582 7552 1014
rect 7648 582 7884 1014
rect 7980 582 8216 1014
rect 8312 582 8548 1014
rect 8644 582 8880 1014
rect 8976 582 9212 1014
rect 9308 582 9544 1014
rect 9640 582 9876 1014
rect 9972 582 10208 1014
rect 10304 582 10540 1014
rect 10636 582 10872 1014
rect 10968 582 11204 1014
rect 11300 582 11536 1014
rect 11632 582 11868 1014
rect 11964 582 12200 1014
rect 12296 582 12532 1014
rect 12628 582 12864 1014
rect 12960 582 13196 1014
rect 13292 582 13528 1014
rect 60 572 147 582
rect 13853 219 14004 1462
rect 25 144 14004 219
rect 25 68 175 144
rect 13853 68 14004 144
rect 25 16 14004 68
<< via1 >>
rect 415 21221 423 25184
rect 423 21221 458 25184
rect 458 21221 467 25184
rect 10008 21202 10060 25165
rect 66 16924 141 20888
rect 507 11356 580 15488
rect 10311 21202 10363 25165
rect 13596 21207 13648 25170
rect 13893 16918 13967 20884
rect 9668 15278 9914 15360
rect 9977 14828 10045 15046
rect 6975 14117 7481 14198
rect 6902 13432 6967 13616
rect 6656 13168 6715 13326
rect 7031 13260 7090 13418
rect 7581 14199 7744 14215
rect 7581 13979 7613 14199
rect 7613 13979 7688 14199
rect 7688 13979 7744 14199
rect 7193 13103 7350 13264
rect 7291 12856 7348 13023
rect 8212 14200 8375 14210
rect 8212 13974 8254 14200
rect 8254 13974 8329 14200
rect 8329 13974 8375 14200
rect 8815 14199 8978 14202
rect 8815 13972 8855 14199
rect 8855 13972 8930 14199
rect 8930 13972 8978 14199
rect 8815 13966 8978 13972
rect 10003 14467 10071 14644
rect 10546 15492 11992 15650
rect 9639 14197 9802 14204
rect 9639 13970 9683 14197
rect 9683 13970 9758 14197
rect 9758 13970 9802 14197
rect 9639 13968 9802 13970
rect 7589 13366 7775 13424
rect 9047 13329 9270 13392
rect 9515 13327 9738 13390
rect 10389 14438 10457 14615
rect 10064 13596 10139 13868
rect 9522 12864 9579 13031
rect 8962 12358 9033 12535
rect 6894 11899 7913 12003
rect 8147 11903 8313 12073
rect 8541 11907 8707 12077
rect 8963 11907 9034 12084
rect 9294 11895 9460 12065
rect 9800 11929 10000 11997
rect 9607 11384 9678 11561
rect 9802 11269 10002 11337
rect 10513 13461 10695 13659
rect 10518 12844 10697 13036
rect 10177 11815 10248 11992
rect 10187 11428 10258 11605
rect 10232 11266 10432 11334
rect 10554 10833 11980 10994
rect 13382 14948 13547 15118
rect 12461 11864 12576 11918
rect 13590 14466 13649 14523
rect 13140 13752 13375 13910
rect 13098 13438 13188 13490
rect 13600 13447 13652 13499
rect 13475 12979 13529 13034
rect 13412 12575 13577 12745
rect 368 5766 420 9742
rect 13614 5764 13666 9740
rect 67 1459 142 5440
rect 13894 1462 13967 5428
<< metal2 >>
rect 415 25193 467 25194
rect 0 25184 14034 25193
rect 0 21221 415 25184
rect 467 25170 14034 25184
rect 467 25165 13596 25170
rect 467 21221 10008 25165
rect 0 21202 10008 21221
rect 10060 21202 10311 25165
rect 10363 21207 13596 25165
rect 13648 21207 14034 25170
rect 10363 21202 14034 21207
rect 0 21193 14034 21202
rect 10008 21192 10060 21193
rect 10311 21192 10363 21193
rect 0 20888 14034 20908
rect 0 16924 66 20888
rect 141 20884 14034 20888
rect 141 16924 13893 20884
rect 0 16918 13893 16924
rect 13967 16918 14034 20884
rect 0 16908 14034 16918
rect 423 15488 627 15616
rect 423 11356 507 15488
rect 580 15027 627 15488
rect 580 11515 6203 15027
rect 6658 14324 7864 16908
rect 8835 15715 10041 16908
rect 8835 15360 9914 15715
rect 8835 15278 9668 15360
rect 8835 14324 9914 15278
rect 10514 15650 12005 16086
rect 10514 15492 10546 15650
rect 11992 15492 12005 15650
rect 10514 15480 12005 15492
rect 9977 15046 10045 15056
rect 10514 15046 10710 15480
rect 10045 14829 10710 15046
rect 13102 15118 14034 15134
rect 13102 14948 13382 15118
rect 13547 14948 14034 15118
rect 13102 14934 14034 14948
rect 9977 14818 10045 14828
rect 9993 14467 10003 14644
rect 10071 14547 10081 14644
rect 10389 14615 10457 14625
rect 10071 14467 10389 14547
rect 9993 14460 10389 14467
rect 9993 14457 10138 14460
rect 6658 14215 9914 14324
rect 6658 14198 7581 14215
rect 6658 14117 6975 14198
rect 7481 14117 7581 14198
rect 6658 13979 7581 14117
rect 7744 14210 9914 14215
rect 7744 13979 8212 14210
rect 6658 13974 8212 13979
rect 8375 14204 9914 14210
rect 8375 14202 9639 14204
rect 8375 13974 8815 14202
rect 6658 13966 8815 13974
rect 8978 13968 9639 14202
rect 9802 13968 9914 14204
rect 8978 13966 9914 13968
rect 6658 13877 9914 13966
rect 10064 13874 10138 14457
rect 10389 14428 10457 14438
rect 10064 13868 10139 13874
rect 6902 13616 6967 13626
rect 10514 13669 10710 14829
rect 13020 14704 13529 14758
rect 13114 13926 13395 13928
rect 13114 13910 13411 13926
rect 13114 13752 13140 13910
rect 13375 13752 13411 13910
rect 13114 13730 13411 13752
rect 10064 13586 10139 13596
rect 10513 13659 10710 13669
rect 6967 13499 9856 13551
rect 6902 13422 6967 13432
rect 7031 13418 7090 13428
rect 6656 13326 6715 13336
rect 6715 13277 7031 13322
rect 7589 13424 7775 13434
rect 7090 13371 7589 13416
rect 9804 13409 9856 13499
rect 10695 13461 10710 13659
rect 13098 13490 13188 13500
rect 10513 13460 10710 13461
rect 10513 13451 10695 13460
rect 12389 13438 13098 13489
rect 12389 13437 13188 13438
rect 12389 13409 12441 13437
rect 13098 13429 13188 13437
rect 7589 13356 7775 13366
rect 9047 13398 9270 13402
rect 9515 13398 9738 13400
rect 9047 13392 9738 13398
rect 9270 13390 9738 13392
rect 9270 13329 9515 13390
rect 9047 13327 9515 13329
rect 9804 13357 12441 13409
rect 9047 13323 9738 13327
rect 9047 13319 9270 13323
rect 9515 13317 9738 13323
rect 7193 13264 7350 13274
rect 13245 13264 13411 13730
rect 7031 13250 7090 13260
rect 6656 13158 6715 13168
rect 7184 13103 7193 13264
rect 7350 13103 13411 13264
rect 7193 13093 7350 13103
rect 7291 13023 7348 13033
rect 9522 13031 9579 13041
rect 7348 12953 9522 13014
rect 7291 12846 7348 12856
rect 9522 12854 9579 12864
rect 10518 13037 10697 13046
rect 10518 13036 10702 13037
rect 10697 12844 10702 13036
rect 10518 12834 10702 12844
rect 8962 12535 9033 12545
rect 8962 12348 9033 12358
rect 6657 12077 8768 12110
rect 8971 12094 9019 12348
rect 6657 12073 8541 12077
rect 6657 12003 8147 12073
rect 6657 11899 6894 12003
rect 7913 11903 8147 12003
rect 8313 11907 8541 12073
rect 8707 11907 8768 12077
rect 8313 11903 8768 11907
rect 7913 11899 8768 11903
rect 6657 11637 8768 11899
rect 8963 12084 9034 12094
rect 8963 11897 9034 11907
rect 9113 12065 9509 12107
rect 9113 11895 9294 12065
rect 9460 11895 9509 12065
rect 9800 12002 10000 12007
rect 10177 12002 10248 12004
rect 9800 11997 10248 12002
rect 10000 11992 10248 11997
rect 10000 11929 10177 11992
rect 9800 11919 10000 11929
rect 9113 11637 9509 11895
rect 10177 11804 10248 11815
rect 580 11356 627 11515
rect 423 9756 627 11356
rect 6657 11084 9509 11637
rect 10187 11605 10258 11615
rect 9607 11561 9678 11571
rect 9678 11472 10187 11534
rect 10187 11418 10258 11428
rect 9607 11374 9678 11384
rect 9802 11337 10002 11347
rect 10232 11334 10432 11344
rect 10002 11272 10232 11330
rect 9802 11259 10002 11269
rect 10232 11256 10432 11266
rect 6657 9756 7863 11084
rect 8830 10951 9509 11084
rect 10525 11031 10702 12834
rect 13245 12759 13411 13103
rect 13475 13034 13529 14704
rect 13590 14523 13649 14533
rect 13834 14523 14034 14657
rect 13649 14466 14034 14523
rect 13590 14456 13649 14466
rect 13834 14457 14034 14466
rect 13600 13509 13639 14456
rect 13600 13499 13652 13509
rect 13600 13437 13652 13447
rect 13600 13429 13639 13437
rect 13475 12966 13529 12979
rect 13245 12745 13577 12759
rect 13245 12575 13412 12745
rect 13577 12575 14034 12659
rect 13245 12459 14034 12575
rect 13834 12105 14034 12174
rect 13247 12051 14034 12105
rect 13834 11974 14034 12051
rect 12461 11918 12576 11928
rect 12461 11854 12576 11864
rect 10525 10994 12010 11031
rect 8830 9756 10036 10951
rect 10525 10833 10554 10994
rect 11980 10833 12010 10994
rect 10525 9756 12010 10833
rect 0 9742 14034 9756
rect 0 5766 368 9742
rect 420 9740 14034 9742
rect 420 5766 13614 9740
rect 0 5764 13614 5766
rect 13666 5764 14034 9740
rect 0 5756 14034 5764
rect 13614 5754 13666 5756
rect 67 5448 142 5450
rect 0 5440 14034 5448
rect 0 1459 67 5440
rect 142 5428 14034 5440
rect 142 1462 13894 5428
rect 13967 1462 14034 5428
rect 142 1459 14034 1462
rect 0 1448 14034 1459
use sky130_fd_pr__diode_pd2nw_05v5_K4SERG  D1
timestamp 1698702074
transform 1 0 9814 0 1 15473
box -321 -321 321 321
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D2
timestamp 1698702074
transform 1 0 9160 0 1 15470
box -183 -183 183 183
use level_shifter  level_shifter_0
timestamp 1698861938
transform -1 0 13172 0 -1 13219
box -422 -2464 2736 144
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  sky130_fd_pr__diode_pw2nd_05v5_FT76RJ_0
timestamp 1698702074
transform 1 0 13785 0 1 14784
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  sky130_fd_pr__diode_pw2nd_05v5_FT76RJ_1
timestamp 1698702074
transform 1 0 12555 0 1 11309
box -183 -183 183 183
use sky130_fd_pr__pfet_01v8_LGS3BL  sky130_fd_pr__pfet_01v8_LGS3BL_0
timestamp 1698716925
transform -1 0 13823 0 1 14142
box -211 -284 211 284
use level_shifter  x2
timestamp 1698861938
transform -1 0 13172 0 1 13291
box -422 -2464 2736 144
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM1
timestamp 1698788623
transform -1 0 8714 0 1 12953
box -278 -269 278 269
use sky130_fd_pr__pfet_g5v0d10v5_XHZHTH  XM2
timestamp 1698788623
transform -1 0 8990 0 1 13744
box -308 -304 308 304
use sky130_fd_pr__pfet_g5v0d10v5_XHZHTH  XM3
timestamp 1698788623
transform -1 0 8374 0 1 13744
box -308 -304 308 304
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM4
timestamp 1698788623
transform -1 0 8158 0 1 12953
box -278 -269 278 269
use sky130_fd_pr__nfet_01v8_L9WNCD  XM5
timestamp 1698716925
transform -1 0 13410 0 -1 13391
box -211 -229 211 229
use sky130_fd_pr__pfet_g5v0d10v5_XHZHTH  XM9
timestamp 1698788623
transform -1 0 7758 0 1 13744
box -308 -304 308 304
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM10
timestamp 1698788623
transform -1 0 7602 0 1 12953
box -278 -269 278 269
use sky130_fd_pr__pfet_g5v0d10v5_XHZHTH  XM11
timestamp 1698788623
transform -1 0 7142 0 1 13744
box -308 -304 308 304
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM12
timestamp 1698788623
transform -1 0 7046 0 -1 12353
box -278 -269 278 269
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM13
timestamp 1698788623
transform -1 0 7046 0 1 12953
box -278 -269 278 269
use sky130_fd_pr__nfet_01v8_L9KS9E  XM14
timestamp 1698716925
transform -1 0 13823 0 1 13391
box -211 -229 211 229
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM21
timestamp 1698788623
transform -1 0 9826 0 -1 12353
box -278 -269 278 269
use sky130_fd_pr__pfet_g5v0d10v5_XHZHTH  XM22
timestamp 1698788623
transform -1 0 9606 0 1 13744
box -308 -304 308 304
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM23
timestamp 1698788623
transform -1 0 9826 0 1 12953
box -278 -269 278 269
use sky130_fd_pr__pfet_g5v0d10v5_XHZHTH  XM24
timestamp 1698788623
transform -1 0 8990 0 -1 14422
box -308 -304 308 304
use sky130_fd_pr__pfet_g5v0d10v5_XHZHTH  XM25
timestamp 1698788623
transform -1 0 8374 0 -1 14422
box -308 -304 308 304
use sky130_fd_pr__pfet_g5v0d10v5_XHZHTH  XM26
timestamp 1698788623
transform -1 0 7758 0 -1 14422
box -308 -304 308 304
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM27
timestamp 1698788623
transform -1 0 7602 0 -1 12353
box -278 -269 278 269
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM28
timestamp 1698788623
transform -1 0 8158 0 -1 12353
box -278 -269 278 269
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM29
timestamp 1698788623
transform -1 0 8714 0 -1 12353
box -278 -269 278 269
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM30
timestamp 1698788623
transform -1 0 9270 0 -1 12353
box -278 -269 278 269
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM31
timestamp 1698788623
transform -1 0 8716 0 -1 11627
box -278 -269 278 269
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM32
timestamp 1698788623
transform -1 0 8160 0 -1 11627
box -278 -269 278 269
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM33
timestamp 1698788623
transform -1 0 9272 0 -1 11627
box -278 -269 278 269
use sky130_fd_pr__pfet_g5v0d10v5_XHZHTH  XM34
timestamp 1698788623
transform -1 0 9606 0 -1 14422
box -308 -304 308 304
use sky130_fd_pr__nfet_01v8_L78EGD  XM35
timestamp 1698716925
transform -1 0 13823 0 1 12941
box -211 -221 211 221
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM36
timestamp 1698788623
transform -1 0 9270 0 1 12953
box -278 -269 278 269
use sky130_fd_pr__nfet_g5v0d10v5_ZFATWT  XM46
timestamp 1698788623
transform -1 0 9828 0 -1 11627
box -278 -269 278 269
use sky130_fd_pr__res_xhigh_po_0p35_6T4SHR  XR1
timestamp 1698702074
transform 1 0 7019 0 1 5498
box -6675 -5082 6675 5082
use sky130_fd_pr__res_high_po_0p69_7CN4E3  XR2
timestamp 1698702074
transform 1 0 3430 0 1 13264
box -2926 -2482 2926 2482
use sky130_fd_pr__res_xhigh_po_0p35_6T4E5R  XR3
timestamp 1698702074
transform -1 0 5237 0 1 21076
box -4849 -5082 4849 5082
use sky130_fd_pr__res_xhigh_po_0p35_9AHPBN  XR4
timestamp 1698702074
transform -1 0 11979 0 1 21066
box -1695 -5082 1695 5082
use sky130_fd_pr__res_high_po_0p69_CY6CB8  XR8
timestamp 1698702074
transform -1 0 12687 0 -1 13238
box -235 -1582 235 1582
<< labels >>
flabel metal1 0 11009 200 11209 0 FreeSans 800 0 0 0 out
port 1 nsew
flabel metal1 0 26179 200 26379 0 FreeSans 800 0 0 0 in
port 0 nsew
flabel metal1 13834 15297 14034 15497 0 FreeSans 800 0 0 0 dout
port 7 nsew
flabel metal2 13834 14934 14034 15134 0 FreeSans 800 0 0 0 dvss
port 4 nsew
flabel metal2 13834 14457 14034 14657 0 FreeSans 800 0 0 0 ena
port 6 nsew
flabel metal2 13834 12459 14034 12659 0 FreeSans 800 0 0 0 dvdd
port 5 nsew
flabel metal2 13834 11974 14034 12174 0 FreeSans 800 0 0 0 boost
port 8 nsew
flabel metal2 s 0 16908 342 20908 0 FreeSans 1280 90 0 0 avdd
port 2 nsew
flabel metal2 0 5756 342 9756 0 FreeSans 1280 90 0 0 avss
port 3 nsew
flabel metal2 13692 5756 14034 9756 0 FreeSans 1280 90 0 0 avss
port 3 nsew
flabel metal2 0 21193 342 25193 0 FreeSans 1280 90 0 0 avss
port 3 nsew
flabel metal2 13692 21193 14034 25193 0 FreeSans 1280 90 0 0 avss
port 3 nsew
flabel metal2 s 13692 16908 14034 20908 0 FreeSans 1280 90 0 0 avdd
port 2 nsew
flabel metal2 s 0 1448 342 5448 0 FreeSans 1280 90 0 0 avdd
port 2 nsew
flabel metal2 s 13692 1448 14034 5448 0 FreeSans 1280 90 0 0 avdd
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 14034 26558
<< end >>
